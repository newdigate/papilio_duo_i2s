----------------------------------------------------------------------
--                                                                  --
--  THIS VHDL SOURCE CODE IS PROVIDED UNDER THE GNU PUBLIC LICENSE  --
--                                                                  --
----------------------------------------------------------------------
--                                                                  --
--    Filename            : sincos_lut.vhd                          --
--                                                                  --
--    Author              : Simon Doherty                           --
--                          Senior Design Consultant                --
--                          www.zipcores.com                        --
--                                                                  --
--    Date last modified  : 26.05.2008                              --
--                                                                  --
--    Description         : 4096 x 12-bit SIN/COS Look-up table     --
--                                                                  --
----------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity sincos_lut_14addr_16 is

port (

  clk       : in  std_logic;
  addr      : in  std_logic_vector(13 downto 0);
  addr_1    : in  std_logic_vector(13 downto 0);
  sin_out   : out std_logic_vector(15 downto 0);
  sin_out_1 : out std_logic_vector(15 downto 0)
  );
  
end entity;


 architecture rtl of sincos_lut_14addr_16 is


type rom_type is array (0 to 16383) of std_logic_vector (15 downto 0);

constant SIN_ROM : rom_type :=

(
X"0000", X"000d", X"0019", X"0026", X"0032", X"003f", X"004b", X"0058", 
X"0065", X"0071", X"007e", X"008a", X"0097", X"00a3", X"00b0", X"00bc", 
X"00c9", X"00d6", X"00e2", X"00ef", X"00fb", X"0108", X"0114", X"0121", 
X"012e", X"013a", X"0147", X"0153", X"0160", X"016c", X"0179", X"0186", 
X"0192", X"019f", X"01ab", X"01b8", X"01c4", X"01d1", X"01de", X"01ea", 
X"01f7", X"0203", X"0210", X"021c", X"0229", X"0235", X"0242", X"024f", 
X"025b", X"0268", X"0274", X"0281", X"028d", X"029a", X"02a7", X"02b3", 
X"02c0", X"02cc", X"02d9", X"02e5", X"02f2", X"02fe", X"030b", X"0318", 
X"0324", X"0331", X"033d", X"034a", X"0356", X"0363", X"0370", X"037c", 
X"0389", X"0395", X"03a2", X"03ae", X"03bb", X"03c7", X"03d4", X"03e1", 
X"03ed", X"03fa", X"0406", X"0413", X"041f", X"042c", X"0439", X"0445", 
X"0452", X"045e", X"046b", X"0477", X"0484", X"0490", X"049d", X"04aa", 
X"04b6", X"04c3", X"04cf", X"04dc", X"04e8", X"04f5", X"0501", X"050e", 
X"051b", X"0527", X"0534", X"0540", X"054d", X"0559", X"0566", X"0572", 
X"057f", X"058c", X"0598", X"05a5", X"05b1", X"05be", X"05ca", X"05d7", 
X"05e3", X"05f0", X"05fd", X"0609", X"0616", X"0622", X"062f", X"063b", 
X"0648", X"0654", X"0661", X"066e", X"067a", X"0687", X"0693", X"06a0", 
X"06ac", X"06b9", X"06c5", X"06d2", X"06de", X"06eb", X"06f8", X"0704", 
X"0711", X"071d", X"072a", X"0736", X"0743", X"074f", X"075c", X"0768", 
X"0775", X"0782", X"078e", X"079b", X"07a7", X"07b4", X"07c0", X"07cd", 
X"07d9", X"07e6", X"07f2", X"07ff", X"080c", X"0818", X"0825", X"0831", 
X"083e", X"084a", X"0857", X"0863", X"0870", X"087c", X"0889", X"0895", 
X"08a2", X"08af", X"08bb", X"08c8", X"08d4", X"08e1", X"08ed", X"08fa", 
X"0906", X"0913", X"091f", X"092c", X"0938", X"0945", X"0951", X"095e", 
X"096b", X"0977", X"0984", X"0990", X"099d", X"09a9", X"09b6", X"09c2", 
X"09cf", X"09db", X"09e8", X"09f4", X"0a01", X"0a0d", X"0a1a", X"0a27", 
X"0a33", X"0a40", X"0a4c", X"0a59", X"0a65", X"0a72", X"0a7e", X"0a8b", 
X"0a97", X"0aa4", X"0ab0", X"0abd", X"0ac9", X"0ad6", X"0ae2", X"0aef", 
X"0afb", X"0b08", X"0b14", X"0b21", X"0b2d", X"0b3a", X"0b47", X"0b53", 
X"0b60", X"0b6c", X"0b79", X"0b85", X"0b92", X"0b9e", X"0bab", X"0bb7", 
X"0bc4", X"0bd0", X"0bdd", X"0be9", X"0bf6", X"0c02", X"0c0f", X"0c1b", 
X"0c28", X"0c34", X"0c41", X"0c4d", X"0c5a", X"0c66", X"0c73", X"0c7f", 
X"0c8c", X"0c98", X"0ca5", X"0cb1", X"0cbe", X"0cca", X"0cd7", X"0ce3", 
X"0cf0", X"0cfc", X"0d09", X"0d15", X"0d22", X"0d2e", X"0d3b", X"0d47", 
X"0d54", X"0d60", X"0d6d", X"0d79", X"0d86", X"0d92", X"0d9f", X"0dab", 
X"0db8", X"0dc4", X"0dd1", X"0ddd", X"0dea", X"0df6", X"0e03", X"0e0f", 
X"0e1c", X"0e28", X"0e35", X"0e41", X"0e4e", X"0e5a", X"0e67", X"0e73", 
X"0e80", X"0e8c", X"0e99", X"0ea5", X"0eb2", X"0ebe", X"0ecb", X"0ed7", 
X"0ee4", X"0ef0", X"0efc", X"0f09", X"0f15", X"0f22", X"0f2e", X"0f3b", 
X"0f47", X"0f54", X"0f60", X"0f6d", X"0f79", X"0f86", X"0f92", X"0f9f", 
X"0fab", X"0fb8", X"0fc4", X"0fd1", X"0fdd", X"0fea", X"0ff6", X"1002", 
X"100f", X"101b", X"1028", X"1034", X"1041", X"104d", X"105a", X"1066", 
X"1073", X"107f", X"108c", X"1098", X"10a4", X"10b1", X"10bd", X"10ca", 
X"10d6", X"10e3", X"10ef", X"10fc", X"1108", X"1115", X"1121", X"112d", 
X"113a", X"1146", X"1153", X"115f", X"116c", X"1178", X"1185", X"1191", 
X"119e", X"11aa", X"11b6", X"11c3", X"11cf", X"11dc", X"11e8", X"11f5", 
X"1201", X"120e", X"121a", X"1226", X"1233", X"123f", X"124c", X"1258", 
X"1265", X"1271", X"127d", X"128a", X"1296", X"12a3", X"12af", X"12bc", 
X"12c8", X"12d4", X"12e1", X"12ed", X"12fa", X"1306", X"1313", X"131f", 
X"132b", X"1338", X"1344", X"1351", X"135d", X"136a", X"1376", X"1382", 
X"138f", X"139b", X"13a8", X"13b4", X"13c1", X"13cd", X"13d9", X"13e6", 
X"13f2", X"13ff", X"140b", X"1417", X"1424", X"1430", X"143d", X"1449", 
X"1455", X"1462", X"146e", X"147b", X"1487", X"1493", X"14a0", X"14ac", 
X"14b9", X"14c5", X"14d1", X"14de", X"14ea", X"14f7", X"1503", X"150f", 
X"151c", X"1528", X"1535", X"1541", X"154d", X"155a", X"1566", X"1573", 
X"157f", X"158b", X"1598", X"15a4", X"15b1", X"15bd", X"15c9", X"15d6", 
X"15e2", X"15ee", X"15fb", X"1607", X"1614", X"1620", X"162c", X"1639", 
X"1645", X"1651", X"165e", X"166a", X"1677", X"1683", X"168f", X"169c", 
X"16a8", X"16b4", X"16c1", X"16cd", X"16da", X"16e6", X"16f2", X"16ff", 
X"170b", X"1717", X"1724", X"1730", X"173c", X"1749", X"1755", X"1761", 
X"176e", X"177a", X"1787", X"1793", X"179f", X"17ac", X"17b8", X"17c4", 
X"17d1", X"17dd", X"17e9", X"17f6", X"1802", X"180e", X"181b", X"1827", 
X"1833", X"1840", X"184c", X"1858", X"1865", X"1871", X"187d", X"188a", 
X"1896", X"18a2", X"18af", X"18bb", X"18c7", X"18d4", X"18e0", X"18ec", 
X"18f9", X"1905", X"1911", X"191e", X"192a", X"1936", X"1943", X"194f", 
X"195b", X"1968", X"1974", X"1980", X"198d", X"1999", X"19a5", X"19b1", 
X"19be", X"19ca", X"19d6", X"19e3", X"19ef", X"19fb", X"1a08", X"1a14", 
X"1a20", X"1a2d", X"1a39", X"1a45", X"1a51", X"1a5e", X"1a6a", X"1a76", 
X"1a83", X"1a8f", X"1a9b", X"1aa8", X"1ab4", X"1ac0", X"1acc", X"1ad9", 
X"1ae5", X"1af1", X"1afe", X"1b0a", X"1b16", X"1b22", X"1b2f", X"1b3b", 
X"1b47", X"1b53", X"1b60", X"1b6c", X"1b78", X"1b85", X"1b91", X"1b9d", 
X"1ba9", X"1bb6", X"1bc2", X"1bce", X"1bda", X"1be7", X"1bf3", X"1bff", 
X"1c0c", X"1c18", X"1c24", X"1c30", X"1c3d", X"1c49", X"1c55", X"1c61", 
X"1c6e", X"1c7a", X"1c86", X"1c92", X"1c9f", X"1cab", X"1cb7", X"1cc3", 
X"1cd0", X"1cdc", X"1ce8", X"1cf4", X"1d01", X"1d0d", X"1d19", X"1d25", 
X"1d31", X"1d3e", X"1d4a", X"1d56", X"1d62", X"1d6f", X"1d7b", X"1d87", 
X"1d93", X"1da0", X"1dac", X"1db8", X"1dc4", X"1dd0", X"1ddd", X"1de9", 
X"1df5", X"1e01", X"1e0e", X"1e1a", X"1e26", X"1e32", X"1e3e", X"1e4b", 
X"1e57", X"1e63", X"1e6f", X"1e7b", X"1e88", X"1e94", X"1ea0", X"1eac", 
X"1eb8", X"1ec5", X"1ed1", X"1edd", X"1ee9", X"1ef5", X"1f02", X"1f0e", 
X"1f1a", X"1f26", X"1f32", X"1f3f", X"1f4b", X"1f57", X"1f63", X"1f6f", 
X"1f7b", X"1f88", X"1f94", X"1fa0", X"1fac", X"1fb8", X"1fc5", X"1fd1", 
X"1fdd", X"1fe9", X"1ff5", X"2001", X"200e", X"201a", X"2026", X"2032", 
X"203e", X"204a", X"2057", X"2063", X"206f", X"207b", X"2087", X"2093", 
X"209f", X"20ac", X"20b8", X"20c4", X"20d0", X"20dc", X"20e8", X"20f4", 
X"2101", X"210d", X"2119", X"2125", X"2131", X"213d", X"2149", X"2156", 
X"2162", X"216e", X"217a", X"2186", X"2192", X"219e", X"21aa", X"21b7", 
X"21c3", X"21cf", X"21db", X"21e7", X"21f3", X"21ff", X"220b", X"2218", 
X"2224", X"2230", X"223c", X"2248", X"2254", X"2260", X"226c", X"2278", 
X"2284", X"2291", X"229d", X"22a9", X"22b5", X"22c1", X"22cd", X"22d9", 
X"22e5", X"22f1", X"22fd", X"230a", X"2316", X"2322", X"232e", X"233a", 
X"2346", X"2352", X"235e", X"236a", X"2376", X"2382", X"238e", X"239a", 
X"23a7", X"23b3", X"23bf", X"23cb", X"23d7", X"23e3", X"23ef", X"23fb", 
X"2407", X"2413", X"241f", X"242b", X"2437", X"2443", X"244f", X"245b", 
X"2467", X"2474", X"2480", X"248c", X"2498", X"24a4", X"24b0", X"24bc", 
X"24c8", X"24d4", X"24e0", X"24ec", X"24f8", X"2504", X"2510", X"251c", 
X"2528", X"2534", X"2540", X"254c", X"2558", X"2564", X"2570", X"257c", 
X"2588", X"2594", X"25a0", X"25ac", X"25b8", X"25c4", X"25d0", X"25dc", 
X"25e8", X"25f4", X"2600", X"260c", X"2618", X"2624", X"2630", X"263c", 
X"2648", X"2654", X"2660", X"266c", X"2678", X"2684", X"2690", X"269c", 
X"26a8", X"26b4", X"26c0", X"26cc", X"26d8", X"26e4", X"26f0", X"26fc", 
X"2708", X"2714", X"2720", X"272c", X"2738", X"2744", X"2750", X"275c", 
X"2768", X"2774", X"2780", X"278b", X"2797", X"27a3", X"27af", X"27bb", 
X"27c7", X"27d3", X"27df", X"27eb", X"27f7", X"2803", X"280f", X"281b", 
X"2827", X"2833", X"283f", X"284b", X"2856", X"2862", X"286e", X"287a", 
X"2886", X"2892", X"289e", X"28aa", X"28b6", X"28c2", X"28ce", X"28da", 
X"28e5", X"28f1", X"28fd", X"2909", X"2915", X"2921", X"292d", X"2939", 
X"2945", X"2951", X"295c", X"2968", X"2974", X"2980", X"298c", X"2998", 
X"29a4", X"29b0", X"29bc", X"29c7", X"29d3", X"29df", X"29eb", X"29f7", 
X"2a03", X"2a0f", X"2a1b", X"2a26", X"2a32", X"2a3e", X"2a4a", X"2a56", 
X"2a62", X"2a6e", X"2a79", X"2a85", X"2a91", X"2a9d", X"2aa9", X"2ab5", 
X"2ac1", X"2acc", X"2ad8", X"2ae4", X"2af0", X"2afc", X"2b08", X"2b13", 
X"2b1f", X"2b2b", X"2b37", X"2b43", X"2b4f", X"2b5a", X"2b66", X"2b72", 
X"2b7e", X"2b8a", X"2b95", X"2ba1", X"2bad", X"2bb9", X"2bc5", X"2bd0", 
X"2bdc", X"2be8", X"2bf4", X"2c00", X"2c0c", X"2c17", X"2c23", X"2c2f", 
X"2c3b", X"2c46", X"2c52", X"2c5e", X"2c6a", X"2c76", X"2c81", X"2c8d", 
X"2c99", X"2ca5", X"2cb1", X"2cbc", X"2cc8", X"2cd4", X"2ce0", X"2ceb", 
X"2cf7", X"2d03", X"2d0f", X"2d1a", X"2d26", X"2d32", X"2d3e", X"2d49", 
X"2d55", X"2d61", X"2d6d", X"2d78", X"2d84", X"2d90", X"2d9c", X"2da7", 
X"2db3", X"2dbf", X"2dcb", X"2dd6", X"2de2", X"2dee", X"2dfa", X"2e05", 
X"2e11", X"2e1d", X"2e28", X"2e34", X"2e40", X"2e4c", X"2e57", X"2e63", 
X"2e6f", X"2e7a", X"2e86", X"2e92", X"2e9e", X"2ea9", X"2eb5", X"2ec1", 
X"2ecc", X"2ed8", X"2ee4", X"2eef", X"2efb", X"2f07", X"2f13", X"2f1e", 
X"2f2a", X"2f36", X"2f41", X"2f4d", X"2f59", X"2f64", X"2f70", X"2f7c", 
X"2f87", X"2f93", X"2f9f", X"2faa", X"2fb6", X"2fc2", X"2fcd", X"2fd9", 
X"2fe5", X"2ff0", X"2ffc", X"3008", X"3013", X"301f", X"302a", X"3036", 
X"3042", X"304d", X"3059", X"3065", X"3070", X"307c", X"3088", X"3093", 
X"309f", X"30aa", X"30b6", X"30c2", X"30cd", X"30d9", X"30e5", X"30f0", 
X"30fc", X"3107", X"3113", X"311f", X"312a", X"3136", X"3141", X"314d", 
X"3159", X"3164", X"3170", X"317b", X"3187", X"3193", X"319e", X"31aa", 
X"31b5", X"31c1", X"31cc", X"31d8", X"31e4", X"31ef", X"31fb", X"3206", 
X"3212", X"321d", X"3229", X"3235", X"3240", X"324c", X"3257", X"3263", 
X"326e", X"327a", X"3285", X"3291", X"329d", X"32a8", X"32b4", X"32bf", 
X"32cb", X"32d6", X"32e2", X"32ed", X"32f9", X"3304", X"3310", X"331b", 
X"3327", X"3332", X"333e", X"3349", X"3355", X"3360", X"336c", X"3377", 
X"3383", X"338e", X"339a", X"33a5", X"33b1", X"33bc", X"33c8", X"33d3", 
X"33df", X"33ea", X"33f6", X"3401", X"340d", X"3418", X"3424", X"342f", 
X"343b", X"3446", X"3452", X"345d", X"3469", X"3474", X"3480", X"348b", 
X"3497", X"34a2", X"34ad", X"34b9", X"34c4", X"34d0", X"34db", X"34e7", 
X"34f2", X"34fe", X"3509", X"3514", X"3520", X"352b", X"3537", X"3542", 
X"354e", X"3559", X"3564", X"3570", X"357b", X"3587", X"3592", X"359d", 
X"35a9", X"35b4", X"35c0", X"35cb", X"35d7", X"35e2", X"35ed", X"35f9", 
X"3604", X"360f", X"361b", X"3626", X"3632", X"363d", X"3648", X"3654", 
X"365f", X"366b", X"3676", X"3681", X"368d", X"3698", X"36a3", X"36af", 
X"36ba", X"36c5", X"36d1", X"36dc", X"36e8", X"36f3", X"36fe", X"370a", 
X"3715", X"3720", X"372c", X"3737", X"3742", X"374e", X"3759", X"3764", 
X"3770", X"377b", X"3786", X"3792", X"379d", X"37a8", X"37b4", X"37bf", 
X"37ca", X"37d5", X"37e1", X"37ec", X"37f7", X"3803", X"380e", X"3819", 
X"3825", X"3830", X"383b", X"3846", X"3852", X"385d", X"3868", X"3874", 
X"387f", X"388a", X"3895", X"38a1", X"38ac", X"38b7", X"38c2", X"38ce", 
X"38d9", X"38e4", X"38f0", X"38fb", X"3906", X"3911", X"391d", X"3928", 
X"3933", X"393e", X"3949", X"3955", X"3960", X"396b", X"3976", X"3982", 
X"398d", X"3998", X"39a3", X"39af", X"39ba", X"39c5", X"39d0", X"39db", 
X"39e7", X"39f2", X"39fd", X"3a08", X"3a13", X"3a1f", X"3a2a", X"3a35", 
X"3a40", X"3a4b", X"3a57", X"3a62", X"3a6d", X"3a78", X"3a83", X"3a8e", 
X"3a9a", X"3aa5", X"3ab0", X"3abb", X"3ac6", X"3ad1", X"3add", X"3ae8", 
X"3af3", X"3afe", X"3b09", X"3b14", X"3b20", X"3b2b", X"3b36", X"3b41", 
X"3b4c", X"3b57", X"3b62", X"3b6d", X"3b79", X"3b84", X"3b8f", X"3b9a", 
X"3ba5", X"3bb0", X"3bbb", X"3bc6", X"3bd2", X"3bdd", X"3be8", X"3bf3", 
X"3bfe", X"3c09", X"3c14", X"3c1f", X"3c2a", X"3c35", X"3c41", X"3c4c", 
X"3c57", X"3c62", X"3c6d", X"3c78", X"3c83", X"3c8e", X"3c99", X"3ca4", 
X"3caf", X"3cba", X"3cc5", X"3cd0", X"3cdc", X"3ce7", X"3cf2", X"3cfd", 
X"3d08", X"3d13", X"3d1e", X"3d29", X"3d34", X"3d3f", X"3d4a", X"3d55", 
X"3d60", X"3d6b", X"3d76", X"3d81", X"3d8c", X"3d97", X"3da2", X"3dad", 
X"3db8", X"3dc3", X"3dce", X"3dd9", X"3de4", X"3def", X"3dfa", X"3e05", 
X"3e10", X"3e1b", X"3e26", X"3e31", X"3e3c", X"3e47", X"3e52", X"3e5d", 
X"3e68", X"3e73", X"3e7e", X"3e89", X"3e94", X"3e9f", X"3eaa", X"3eb5", 
X"3ec0", X"3ecb", X"3ed6", X"3ee1", X"3eec", X"3ef6", X"3f01", X"3f0c", 
X"3f17", X"3f22", X"3f2d", X"3f38", X"3f43", X"3f4e", X"3f59", X"3f64", 
X"3f6f", X"3f7a", X"3f85", X"3f8f", X"3f9a", X"3fa5", X"3fb0", X"3fbb", 
X"3fc6", X"3fd1", X"3fdc", X"3fe7", X"3ff1", X"3ffc", X"4007", X"4012", 
X"401d", X"4028", X"4033", X"403e", X"4048", X"4053", X"405e", X"4069", 
X"4074", X"407f", X"408a", X"4095", X"409f", X"40aa", X"40b5", X"40c0", 
X"40cb", X"40d6", X"40e0", X"40eb", X"40f6", X"4101", X"410c", X"4117", 
X"4121", X"412c", X"4137", X"4142", X"414d", X"4157", X"4162", X"416d", 
X"4178", X"4183", X"418d", X"4198", X"41a3", X"41ae", X"41b9", X"41c3", 
X"41ce", X"41d9", X"41e4", X"41ee", X"41f9", X"4204", X"420f", X"421a", 
X"4224", X"422f", X"423a", X"4245", X"424f", X"425a", X"4265", X"4270", 
X"427a", X"4285", X"4290", X"429a", X"42a5", X"42b0", X"42bb", X"42c5", 
X"42d0", X"42db", X"42e6", X"42f0", X"42fb", X"4306", X"4310", X"431b", 
X"4326", X"4330", X"433b", X"4346", X"4351", X"435b", X"4366", X"4371", 
X"437b", X"4386", X"4391", X"439b", X"43a6", X"43b1", X"43bb", X"43c6", 
X"43d1", X"43db", X"43e6", X"43f1", X"43fb", X"4406", X"4411", X"441b", 
X"4426", X"4430", X"443b", X"4446", X"4450", X"445b", X"4466", X"4470", 
X"447b", X"4485", X"4490", X"449b", X"44a5", X"44b0", X"44ba", X"44c5", 
X"44d0", X"44da", X"44e5", X"44ef", X"44fa", X"4505", X"450f", X"451a", 
X"4524", X"452f", X"4539", X"4544", X"454f", X"4559", X"4564", X"456e", 
X"4579", X"4583", X"458e", X"4599", X"45a3", X"45ae", X"45b8", X"45c3", 
X"45cd", X"45d8", X"45e2", X"45ed", X"45f7", X"4602", X"460c", X"4617", 
X"4621", X"462c", X"4636", X"4641", X"464b", X"4656", X"4660", X"466b", 
X"4675", X"4680", X"468a", X"4695", X"469f", X"46aa", X"46b4", X"46bf", 
X"46c9", X"46d4", X"46de", X"46e9", X"46f3", X"46fe", X"4708", X"4712", 
X"471d", X"4727", X"4732", X"473c", X"4747", X"4751", X"475c", X"4766", 
X"4770", X"477b", X"4785", X"4790", X"479a", X"47a5", X"47af", X"47b9", 
X"47c4", X"47ce", X"47d9", X"47e3", X"47ed", X"47f8", X"4802", X"480d", 
X"4817", X"4821", X"482c", X"4836", X"4840", X"484b", X"4855", X"4860", 
X"486a", X"4874", X"487f", X"4889", X"4893", X"489e", X"48a8", X"48b2", 
X"48bd", X"48c7", X"48d1", X"48dc", X"48e6", X"48f0", X"48fb", X"4905", 
X"490f", X"491a", X"4924", X"492e", X"4939", X"4943", X"494d", X"4958", 
X"4962", X"496c", X"4976", X"4981", X"498b", X"4995", X"49a0", X"49aa", 
X"49b4", X"49be", X"49c9", X"49d3", X"49dd", X"49e7", X"49f2", X"49fc", 
X"4a06", X"4a10", X"4a1b", X"4a25", X"4a2f", X"4a39", X"4a44", X"4a4e", 
X"4a58", X"4a62", X"4a6d", X"4a77", X"4a81", X"4a8b", X"4a95", X"4aa0", 
X"4aaa", X"4ab4", X"4abe", X"4ac8", X"4ad3", X"4add", X"4ae7", X"4af1", 
X"4afb", X"4b06", X"4b10", X"4b1a", X"4b24", X"4b2e", X"4b38", X"4b43", 
X"4b4d", X"4b57", X"4b61", X"4b6b", X"4b75", X"4b80", X"4b8a", X"4b94", 
X"4b9e", X"4ba8", X"4bb2", X"4bbc", X"4bc7", X"4bd1", X"4bdb", X"4be5", 
X"4bef", X"4bf9", X"4c03", X"4c0d", X"4c17", X"4c22", X"4c2c", X"4c36", 
X"4c40", X"4c4a", X"4c54", X"4c5e", X"4c68", X"4c72", X"4c7c", X"4c86", 
X"4c91", X"4c9b", X"4ca5", X"4caf", X"4cb9", X"4cc3", X"4ccd", X"4cd7", 
X"4ce1", X"4ceb", X"4cf5", X"4cff", X"4d09", X"4d13", X"4d1d", X"4d27", 
X"4d31", X"4d3b", X"4d45", X"4d4f", X"4d59", X"4d63", X"4d6d", X"4d77", 
X"4d81", X"4d8b", X"4d95", X"4d9f", X"4da9", X"4db3", X"4dbd", X"4dc7", 
X"4dd1", X"4ddb", X"4de5", X"4def", X"4df9", X"4e03", X"4e0d", X"4e17", 
X"4e21", X"4e2b", X"4e35", X"4e3f", X"4e49", X"4e53", X"4e5d", X"4e67", 
X"4e71", X"4e7a", X"4e84", X"4e8e", X"4e98", X"4ea2", X"4eac", X"4eb6", 
X"4ec0", X"4eca", X"4ed4", X"4ede", X"4ee8", X"4ef1", X"4efb", X"4f05", 
X"4f0f", X"4f19", X"4f23", X"4f2d", X"4f37", X"4f40", X"4f4a", X"4f54", 
X"4f5e", X"4f68", X"4f72", X"4f7c", X"4f85", X"4f8f", X"4f99", X"4fa3", 
X"4fad", X"4fb7", X"4fc0", X"4fca", X"4fd4", X"4fde", X"4fe8", X"4ff2", 
X"4ffb", X"5005", X"500f", X"5019", X"5023", X"502c", X"5036", X"5040", 
X"504a", X"5054", X"505d", X"5067", X"5071", X"507b", X"5084", X"508e", 
X"5098", X"50a2", X"50ac", X"50b5", X"50bf", X"50c9", X"50d3", X"50dc", 
X"50e6", X"50f0", X"50f9", X"5103", X"510d", X"5117", X"5120", X"512a", 
X"5134", X"513e", X"5147", X"5151", X"515b", X"5164", X"516e", X"5178", 
X"5181", X"518b", X"5195", X"519e", X"51a8", X"51b2", X"51bb", X"51c5", 
X"51cf", X"51d8", X"51e2", X"51ec", X"51f5", X"51ff", X"5209", X"5212", 
X"521c", X"5226", X"522f", X"5239", X"5243", X"524c", X"5256", X"525f", 
X"5269", X"5273", X"527c", X"5286", X"5290", X"5299", X"52a3", X"52ac", 
X"52b6", X"52bf", X"52c9", X"52d3", X"52dc", X"52e6", X"52ef", X"52f9", 
X"5303", X"530c", X"5316", X"531f", X"5329", X"5332", X"533c", X"5345", 
X"534f", X"5358", X"5362", X"536c", X"5375", X"537f", X"5388", X"5392", 
X"539b", X"53a5", X"53ae", X"53b8", X"53c1", X"53cb", X"53d4", X"53de", 
X"53e7", X"53f1", X"53fa", X"5404", X"540d", X"5417", X"5420", X"542a", 
X"5433", X"543c", X"5446", X"544f", X"5459", X"5462", X"546c", X"5475", 
X"547f", X"5488", X"5491", X"549b", X"54a4", X"54ae", X"54b7", X"54c1", 
X"54ca", X"54d3", X"54dd", X"54e6", X"54f0", X"54f9", X"5502", X"550c", 
X"5515", X"551f", X"5528", X"5531", X"553b", X"5544", X"554e", X"5557", 
X"5560", X"556a", X"5573", X"557c", X"5586", X"558f", X"5598", X"55a2", 
X"55ab", X"55b4", X"55be", X"55c7", X"55d0", X"55da", X"55e3", X"55ec", 
X"55f6", X"55ff", X"5608", X"5612", X"561b", X"5624", X"562d", X"5637", 
X"5640", X"5649", X"5653", X"565c", X"5665", X"566e", X"5678", X"5681", 
X"568a", X"5693", X"569d", X"56a6", X"56af", X"56b8", X"56c2", X"56cb", 
X"56d4", X"56dd", X"56e7", X"56f0", X"56f9", X"5702", X"570c", X"5715", 
X"571e", X"5727", X"5730", X"573a", X"5743", X"574c", X"5755", X"575e", 
X"5767", X"5771", X"577a", X"5783", X"578c", X"5795", X"579f", X"57a8", 
X"57b1", X"57ba", X"57c3", X"57cc", X"57d5", X"57df", X"57e8", X"57f1", 
X"57fa", X"5803", X"580c", X"5815", X"581e", X"5828", X"5831", X"583a", 
X"5843", X"584c", X"5855", X"585e", X"5867", X"5870", X"5879", X"5882", 
X"588c", X"5895", X"589e", X"58a7", X"58b0", X"58b9", X"58c2", X"58cb", 
X"58d4", X"58dd", X"58e6", X"58ef", X"58f8", X"5901", X"590a", X"5913", 
X"591c", X"5925", X"592e", X"5937", X"5940", X"5949", X"5952", X"595b", 
X"5964", X"596d", X"5976", X"597f", X"5988", X"5991", X"599a", X"59a3", 
X"59ac", X"59b5", X"59be", X"59c7", X"59d0", X"59d9", X"59e2", X"59eb", 
X"59f4", X"59fd", X"5a06", X"5a0f", X"5a18", X"5a21", X"5a29", X"5a32", 
X"5a3b", X"5a44", X"5a4d", X"5a56", X"5a5f", X"5a68", X"5a71", X"5a7a", 
X"5a82", X"5a8b", X"5a94", X"5a9d", X"5aa6", X"5aaf", X"5ab8", X"5ac1", 
X"5ac9", X"5ad2", X"5adb", X"5ae4", X"5aed", X"5af6", X"5aff", X"5b07", 
X"5b10", X"5b19", X"5b22", X"5b2b", X"5b34", X"5b3c", X"5b45", X"5b4e", 
X"5b57", X"5b60", X"5b68", X"5b71", X"5b7a", X"5b83", X"5b8c", X"5b94", 
X"5b9d", X"5ba6", X"5baf", X"5bb7", X"5bc0", X"5bc9", X"5bd2", X"5bda", 
X"5be3", X"5bec", X"5bf5", X"5bfd", X"5c06", X"5c0f", X"5c18", X"5c20", 
X"5c29", X"5c32", X"5c3a", X"5c43", X"5c4c", X"5c55", X"5c5d", X"5c66", 
X"5c6f", X"5c77", X"5c80", X"5c89", X"5c91", X"5c9a", X"5ca3", X"5cab", 
X"5cb4", X"5cbd", X"5cc5", X"5cce", X"5cd7", X"5cdf", X"5ce8", X"5cf1", 
X"5cf9", X"5d02", X"5d0b", X"5d13", X"5d1c", X"5d24", X"5d2d", X"5d36", 
X"5d3e", X"5d47", X"5d50", X"5d58", X"5d61", X"5d69", X"5d72", X"5d7a", 
X"5d83", X"5d8c", X"5d94", X"5d9d", X"5da5", X"5dae", X"5db7", X"5dbf", 
X"5dc8", X"5dd0", X"5dd9", X"5de1", X"5dea", X"5df2", X"5dfb", X"5e03", 
X"5e0c", X"5e14", X"5e1d", X"5e25", X"5e2e", X"5e37", X"5e3f", X"5e48", 
X"5e50", X"5e58", X"5e61", X"5e69", X"5e72", X"5e7a", X"5e83", X"5e8b", 
X"5e94", X"5e9c", X"5ea5", X"5ead", X"5eb6", X"5ebe", X"5ec7", X"5ecf", 
X"5ed7", X"5ee0", X"5ee8", X"5ef1", X"5ef9", X"5f02", X"5f0a", X"5f12", 
X"5f1b", X"5f23", X"5f2c", X"5f34", X"5f3c", X"5f45", X"5f4d", X"5f56", 
X"5f5e", X"5f66", X"5f6f", X"5f77", X"5f80", X"5f88", X"5f90", X"5f99", 
X"5fa1", X"5fa9", X"5fb2", X"5fba", X"5fc2", X"5fcb", X"5fd3", X"5fdb", 
X"5fe4", X"5fec", X"5ff4", X"5ffd", X"6005", X"600d", X"6016", X"601e", 
X"6026", X"602e", X"6037", X"603f", X"6047", X"6050", X"6058", X"6060", 
X"6068", X"6071", X"6079", X"6081", X"6089", X"6092", X"609a", X"60a2", 
X"60aa", X"60b3", X"60bb", X"60c3", X"60cb", X"60d4", X"60dc", X"60e4", 
X"60ec", X"60f4", X"60fd", X"6105", X"610d", X"6115", X"611d", X"6126", 
X"612e", X"6136", X"613e", X"6146", X"614e", X"6157", X"615f", X"6167", 
X"616f", X"6177", X"617f", X"6188", X"6190", X"6198", X"61a0", X"61a8", 
X"61b0", X"61b8", X"61c0", X"61c9", X"61d1", X"61d9", X"61e1", X"61e9", 
X"61f1", X"61f9", X"6201", X"6209", X"6211", X"6219", X"6221", X"622a", 
X"6232", X"623a", X"6242", X"624a", X"6252", X"625a", X"6262", X"626a", 
X"6272", X"627a", X"6282", X"628a", X"6292", X"629a", X"62a2", X"62aa", 
X"62b2", X"62ba", X"62c2", X"62ca", X"62d2", X"62da", X"62e2", X"62ea", 
X"62f2", X"62fa", X"6302", X"630a", X"6312", X"631a", X"6322", X"632a", 
X"6332", X"633a", X"6342", X"6349", X"6351", X"6359", X"6361", X"6369", 
X"6371", X"6379", X"6381", X"6389", X"6391", X"6399", X"63a0", X"63a8", 
X"63b0", X"63b8", X"63c0", X"63c8", X"63d0", X"63d8", X"63df", X"63e7", 
X"63ef", X"63f7", X"63ff", X"6407", X"640f", X"6416", X"641e", X"6426", 
X"642e", X"6436", X"643e", X"6445", X"644d", X"6455", X"645d", X"6465", 
X"646c", X"6474", X"647c", X"6484", X"648b", X"6493", X"649b", X"64a3", 
X"64ab", X"64b2", X"64ba", X"64c2", X"64ca", X"64d1", X"64d9", X"64e1", 
X"64e9", X"64f0", X"64f8", X"6500", X"6507", X"650f", X"6517", X"651f", 
X"6526", X"652e", X"6536", X"653d", X"6545", X"654d", X"6554", X"655c", 
X"6564", X"656b", X"6573", X"657b", X"6582", X"658a", X"6592", X"6599", 
X"65a1", X"65a9", X"65b0", X"65b8", X"65c0", X"65c7", X"65cf", X"65d6", 
X"65de", X"65e6", X"65ed", X"65f5", X"65fc", X"6604", X"660c", X"6613", 
X"661b", X"6622", X"662a", X"6631", X"6639", X"6641", X"6648", X"6650", 
X"6657", X"665f", X"6666", X"666e", X"6675", X"667d", X"6684", X"668c", 
X"6693", X"669b", X"66a3", X"66aa", X"66b2", X"66b9", X"66c1", X"66c8", 
X"66d0", X"66d7", X"66de", X"66e6", X"66ed", X"66f5", X"66fc", X"6704", 
X"670b", X"6713", X"671a", X"6722", X"6729", X"6730", X"6738", X"673f", 
X"6747", X"674e", X"6756", X"675d", X"6764", X"676c", X"6773", X"677b", 
X"6782", X"6789", X"6791", X"6798", X"67a0", X"67a7", X"67ae", X"67b6", 
X"67bd", X"67c4", X"67cc", X"67d3", X"67da", X"67e2", X"67e9", X"67f0", 
X"67f8", X"67ff", X"6806", X"680e", X"6815", X"681c", X"6824", X"682b", 
X"6832", X"683a", X"6841", X"6848", X"6850", X"6857", X"685e", X"6865", 
X"686d", X"6874", X"687b", X"6882", X"688a", X"6891", X"6898", X"689f", 
X"68a7", X"68ae", X"68b5", X"68bc", X"68c4", X"68cb", X"68d2", X"68d9", 
X"68e0", X"68e8", X"68ef", X"68f6", X"68fd", X"6904", X"690c", X"6913", 
X"691a", X"6921", X"6928", X"692f", X"6937", X"693e", X"6945", X"694c", 
X"6953", X"695a", X"6961", X"6969", X"6970", X"6977", X"697e", X"6985", 
X"698c", X"6993", X"699a", X"69a1", X"69a9", X"69b0", X"69b7", X"69be", 
X"69c5", X"69cc", X"69d3", X"69da", X"69e1", X"69e8", X"69ef", X"69f6", 
X"69fd", X"6a04", X"6a0b", X"6a12", X"6a1a", X"6a21", X"6a28", X"6a2f", 
X"6a36", X"6a3d", X"6a44", X"6a4b", X"6a52", X"6a59", X"6a60", X"6a67", 
X"6a6e", X"6a75", X"6a7c", X"6a83", X"6a89", X"6a90", X"6a97", X"6a9e", 
X"6aa5", X"6aac", X"6ab3", X"6aba", X"6ac1", X"6ac8", X"6acf", X"6ad6", 
X"6add", X"6ae4", X"6aeb", X"6af2", X"6af8", X"6aff", X"6b06", X"6b0d", 
X"6b14", X"6b1b", X"6b22", X"6b29", X"6b30", X"6b36", X"6b3d", X"6b44", 
X"6b4b", X"6b52", X"6b59", X"6b5f", X"6b66", X"6b6d", X"6b74", X"6b7b", 
X"6b82", X"6b88", X"6b8f", X"6b96", X"6b9d", X"6ba4", X"6baa", X"6bb1", 
X"6bb8", X"6bbf", X"6bc6", X"6bcc", X"6bd3", X"6bda", X"6be1", X"6be7", 
X"6bee", X"6bf5", X"6bfc", X"6c02", X"6c09", X"6c10", X"6c17", X"6c1d", 
X"6c24", X"6c2b", X"6c32", X"6c38", X"6c3f", X"6c46", X"6c4c", X"6c53", 
X"6c5a", X"6c61", X"6c67", X"6c6e", X"6c75", X"6c7b", X"6c82", X"6c89", 
X"6c8f", X"6c96", X"6c9d", X"6ca3", X"6caa", X"6cb0", X"6cb7", X"6cbe", 
X"6cc4", X"6ccb", X"6cd2", X"6cd8", X"6cdf", X"6ce5", X"6cec", X"6cf3", 
X"6cf9", X"6d00", X"6d06", X"6d0d", X"6d14", X"6d1a", X"6d21", X"6d27", 
X"6d2e", X"6d34", X"6d3b", X"6d41", X"6d48", X"6d4f", X"6d55", X"6d5c", 
X"6d62", X"6d69", X"6d6f", X"6d76", X"6d7c", X"6d83", X"6d89", X"6d90", 
X"6d96", X"6d9d", X"6da3", X"6daa", X"6db0", X"6db7", X"6dbd", X"6dc4", 
X"6dca", X"6dd1", X"6dd7", X"6ddd", X"6de4", X"6dea", X"6df1", X"6df7", 
X"6dfe", X"6e04", X"6e0a", X"6e11", X"6e17", X"6e1e", X"6e24", X"6e2a", 
X"6e31", X"6e37", X"6e3e", X"6e44", X"6e4a", X"6e51", X"6e57", X"6e5e", 
X"6e64", X"6e6a", X"6e71", X"6e77", X"6e7d", X"6e84", X"6e8a", X"6e90", 
X"6e97", X"6e9d", X"6ea3", X"6eaa", X"6eb0", X"6eb6", X"6ebd", X"6ec3", 
X"6ec9", X"6ecf", X"6ed6", X"6edc", X"6ee2", X"6ee9", X"6eef", X"6ef5", 
X"6efb", X"6f02", X"6f08", X"6f0e", X"6f14", X"6f1b", X"6f21", X"6f27", 
X"6f2d", X"6f34", X"6f3a", X"6f40", X"6f46", X"6f4c", X"6f53", X"6f59", 
X"6f5f", X"6f65", X"6f6b", X"6f72", X"6f78", X"6f7e", X"6f84", X"6f8a", 
X"6f90", X"6f97", X"6f9d", X"6fa3", X"6fa9", X"6faf", X"6fb5", X"6fbb", 
X"6fc2", X"6fc8", X"6fce", X"6fd4", X"6fda", X"6fe0", X"6fe6", X"6fec", 
X"6ff2", X"6ff9", X"6fff", X"7005", X"700b", X"7011", X"7017", X"701d", 
X"7023", X"7029", X"702f", X"7035", X"703b", X"7041", X"7047", X"704d", 
X"7053", X"7059", X"705f", X"7065", X"706b", X"7071", X"7077", X"707d", 
X"7083", X"7089", X"708f", X"7095", X"709b", X"70a1", X"70a7", X"70ad", 
X"70b3", X"70b9", X"70bf", X"70c5", X"70cb", X"70d1", X"70d7", X"70dd", 
X"70e3", X"70e9", X"70ef", X"70f5", X"70fa", X"7100", X"7106", X"710c", 
X"7112", X"7118", X"711e", X"7124", X"712a", X"712f", X"7135", X"713b", 
X"7141", X"7147", X"714d", X"7153", X"7158", X"715e", X"7164", X"716a", 
X"7170", X"7176", X"717b", X"7181", X"7187", X"718d", X"7193", X"7198", 
X"719e", X"71a4", X"71aa", X"71b0", X"71b5", X"71bb", X"71c1", X"71c7", 
X"71cc", X"71d2", X"71d8", X"71de", X"71e3", X"71e9", X"71ef", X"71f5", 
X"71fa", X"7200", X"7206", X"720b", X"7211", X"7217", X"721c", X"7222", 
X"7228", X"722e", X"7233", X"7239", X"723f", X"7244", X"724a", X"7250", 
X"7255", X"725b", X"7260", X"7266", X"726c", X"7271", X"7277", X"727d", 
X"7282", X"7288", X"728d", X"7293", X"7299", X"729e", X"72a4", X"72a9", 
X"72af", X"72b5", X"72ba", X"72c0", X"72c5", X"72cb", X"72d0", X"72d6", 
X"72dc", X"72e1", X"72e7", X"72ec", X"72f2", X"72f7", X"72fd", X"7302", 
X"7308", X"730d", X"7313", X"7318", X"731e", X"7323", X"7329", X"732e", 
X"7334", X"7339", X"733f", X"7344", X"734a", X"734f", X"7355", X"735a", 
X"735f", X"7365", X"736a", X"7370", X"7375", X"737b", X"7380", X"7385", 
X"738b", X"7390", X"7396", X"739b", X"73a0", X"73a6", X"73ab", X"73b1", 
X"73b6", X"73bb", X"73c1", X"73c6", X"73cb", X"73d1", X"73d6", X"73db", 
X"73e1", X"73e6", X"73eb", X"73f1", X"73f6", X"73fb", X"7401", X"7406", 
X"740b", X"7411", X"7416", X"741b", X"7421", X"7426", X"742b", X"7430", 
X"7436", X"743b", X"7440", X"7445", X"744b", X"7450", X"7455", X"745a", 
X"7460", X"7465", X"746a", X"746f", X"7475", X"747a", X"747f", X"7484", 
X"7489", X"748f", X"7494", X"7499", X"749e", X"74a3", X"74a8", X"74ae", 
X"74b3", X"74b8", X"74bd", X"74c2", X"74c7", X"74cd", X"74d2", X"74d7", 
X"74dc", X"74e1", X"74e6", X"74eb", X"74f0", X"74f6", X"74fb", X"7500", 
X"7505", X"750a", X"750f", X"7514", X"7519", X"751e", X"7523", X"7528", 
X"752d", X"7532", X"7538", X"753d", X"7542", X"7547", X"754c", X"7551", 
X"7556", X"755b", X"7560", X"7565", X"756a", X"756f", X"7574", X"7579", 
X"757e", X"7583", X"7588", X"758d", X"7592", X"7597", X"759c", X"75a1", 
X"75a6", X"75aa", X"75af", X"75b4", X"75b9", X"75be", X"75c3", X"75c8", 
X"75cd", X"75d2", X"75d7", X"75dc", X"75e1", X"75e6", X"75ea", X"75ef", 
X"75f4", X"75f9", X"75fe", X"7603", X"7608", X"760d", X"7611", X"7616", 
X"761b", X"7620", X"7625", X"762a", X"762e", X"7633", X"7638", X"763d", 
X"7642", X"7646", X"764b", X"7650", X"7655", X"765a", X"765e", X"7663", 
X"7668", X"766d", X"7672", X"7676", X"767b", X"7680", X"7685", X"7689", 
X"768e", X"7693", X"7698", X"769c", X"76a1", X"76a6", X"76aa", X"76af", 
X"76b4", X"76b9", X"76bd", X"76c2", X"76c7", X"76cb", X"76d0", X"76d5", 
X"76d9", X"76de", X"76e3", X"76e7", X"76ec", X"76f1", X"76f5", X"76fa", 
X"76fe", X"7703", X"7708", X"770c", X"7711", X"7716", X"771a", X"771f", 
X"7723", X"7728", X"772d", X"7731", X"7736", X"773a", X"773f", X"7743", 
X"7748", X"774d", X"7751", X"7756", X"775a", X"775f", X"7763", X"7768", 
X"776c", X"7771", X"7775", X"777a", X"777e", X"7783", X"7787", X"778c", 
X"7790", X"7795", X"7799", X"779e", X"77a2", X"77a7", X"77ab", X"77b0", 
X"77b4", X"77b9", X"77bd", X"77c1", X"77c6", X"77ca", X"77cf", X"77d3", 
X"77d8", X"77dc", X"77e0", X"77e5", X"77e9", X"77ee", X"77f2", X"77f6", 
X"77fb", X"77ff", X"7803", X"7808", X"780c", X"7811", X"7815", X"7819", 
X"781e", X"7822", X"7826", X"782b", X"782f", X"7833", X"7838", X"783c", 
X"7840", X"7845", X"7849", X"784d", X"7851", X"7856", X"785a", X"785e", 
X"7863", X"7867", X"786b", X"786f", X"7874", X"7878", X"787c", X"7880", 
X"7885", X"7889", X"788d", X"7891", X"7895", X"789a", X"789e", X"78a2", 
X"78a6", X"78aa", X"78af", X"78b3", X"78b7", X"78bb", X"78bf", X"78c4", 
X"78c8", X"78cc", X"78d0", X"78d4", X"78d8", X"78dc", X"78e1", X"78e5", 
X"78e9", X"78ed", X"78f1", X"78f5", X"78f9", X"78fd", X"7901", X"7906", 
X"790a", X"790e", X"7912", X"7916", X"791a", X"791e", X"7922", X"7926", 
X"792a", X"792e", X"7932", X"7936", X"793a", X"793e", X"7942", X"7946", 
X"794a", X"794e", X"7953", X"7957", X"795b", X"795f", X"7962", X"7966", 
X"796a", X"796e", X"7972", X"7976", X"797a", X"797e", X"7982", X"7986", 
X"798a", X"798e", X"7992", X"7996", X"799a", X"799e", X"79a2", X"79a6", 
X"79aa", X"79ad", X"79b1", X"79b5", X"79b9", X"79bd", X"79c1", X"79c5", 
X"79c9", X"79cc", X"79d0", X"79d4", X"79d8", X"79dc", X"79e0", X"79e4", 
X"79e7", X"79eb", X"79ef", X"79f3", X"79f7", X"79fb", X"79fe", X"7a02", 
X"7a06", X"7a0a", X"7a0e", X"7a11", X"7a15", X"7a19", X"7a1d", X"7a20", 
X"7a24", X"7a28", X"7a2c", X"7a2f", X"7a33", X"7a37", X"7a3b", X"7a3e", 
X"7a42", X"7a46", X"7a49", X"7a4d", X"7a51", X"7a55", X"7a58", X"7a5c", 
X"7a60", X"7a63", X"7a67", X"7a6b", X"7a6e", X"7a72", X"7a76", X"7a79", 
X"7a7d", X"7a81", X"7a84", X"7a88", X"7a8c", X"7a8f", X"7a93", X"7a96", 
X"7a9a", X"7a9e", X"7aa1", X"7aa5", X"7aa8", X"7aac", X"7ab0", X"7ab3", 
X"7ab7", X"7aba", X"7abe", X"7ac1", X"7ac5", X"7ac9", X"7acc", X"7ad0", 
X"7ad3", X"7ad7", X"7ada", X"7ade", X"7ae1", X"7ae5", X"7ae8", X"7aec", 
X"7aef", X"7af3", X"7af6", X"7afa", X"7afd", X"7b01", X"7b04", X"7b08", 
X"7b0b", X"7b0f", X"7b12", X"7b16", X"7b19", X"7b1c", X"7b20", X"7b23", 
X"7b27", X"7b2a", X"7b2e", X"7b31", X"7b34", X"7b38", X"7b3b", X"7b3f", 
X"7b42", X"7b45", X"7b49", X"7b4c", X"7b50", X"7b53", X"7b56", X"7b5a", 
X"7b5d", X"7b60", X"7b64", X"7b67", X"7b6a", X"7b6e", X"7b71", X"7b74", 
X"7b78", X"7b7b", X"7b7e", X"7b82", X"7b85", X"7b88", X"7b8b", X"7b8f", 
X"7b92", X"7b95", X"7b99", X"7b9c", X"7b9f", X"7ba2", X"7ba6", X"7ba9", 
X"7bac", X"7baf", X"7bb3", X"7bb6", X"7bb9", X"7bbc", X"7bbf", X"7bc3", 
X"7bc6", X"7bc9", X"7bcc", X"7bcf", X"7bd3", X"7bd6", X"7bd9", X"7bdc", 
X"7bdf", X"7be3", X"7be6", X"7be9", X"7bec", X"7bef", X"7bf2", X"7bf5", 
X"7bf9", X"7bfc", X"7bff", X"7c02", X"7c05", X"7c08", X"7c0b", X"7c0e", 
X"7c11", X"7c14", X"7c18", X"7c1b", X"7c1e", X"7c21", X"7c24", X"7c27", 
X"7c2a", X"7c2d", X"7c30", X"7c33", X"7c36", X"7c39", X"7c3c", X"7c3f", 
X"7c42", X"7c45", X"7c48", X"7c4b", X"7c4e", X"7c51", X"7c54", X"7c57", 
X"7c5a", X"7c5d", X"7c60", X"7c63", X"7c66", X"7c69", X"7c6c", X"7c6f", 
X"7c72", X"7c75", X"7c78", X"7c7b", X"7c7e", X"7c81", X"7c83", X"7c86", 
X"7c89", X"7c8c", X"7c8f", X"7c92", X"7c95", X"7c98", X"7c9b", X"7c9e", 
X"7ca0", X"7ca3", X"7ca6", X"7ca9", X"7cac", X"7caf", X"7cb1", X"7cb4", 
X"7cb7", X"7cba", X"7cbd", X"7cc0", X"7cc2", X"7cc5", X"7cc8", X"7ccb", 
X"7cce", X"7cd0", X"7cd3", X"7cd6", X"7cd9", X"7cdc", X"7cde", X"7ce1", 
X"7ce4", X"7ce7", X"7ce9", X"7cec", X"7cef", X"7cf2", X"7cf4", X"7cf7", 
X"7cfa", X"7cfc", X"7cff", X"7d02", X"7d05", X"7d07", X"7d0a", X"7d0d", 
X"7d0f", X"7d12", X"7d15", X"7d17", X"7d1a", X"7d1d", X"7d1f", X"7d22", 
X"7d25", X"7d27", X"7d2a", X"7d2c", X"7d2f", X"7d32", X"7d34", X"7d37", 
X"7d3a", X"7d3c", X"7d3f", X"7d41", X"7d44", X"7d46", X"7d49", X"7d4c", 
X"7d4e", X"7d51", X"7d53", X"7d56", X"7d58", X"7d5b", X"7d5d", X"7d60", 
X"7d63", X"7d65", X"7d68", X"7d6a", X"7d6d", X"7d6f", X"7d72", X"7d74", 
X"7d77", X"7d79", X"7d7c", X"7d7e", X"7d81", X"7d83", X"7d85", X"7d88", 
X"7d8a", X"7d8d", X"7d8f", X"7d92", X"7d94", X"7d97", X"7d99", X"7d9b", 
X"7d9e", X"7da0", X"7da3", X"7da5", X"7da7", X"7daa", X"7dac", X"7daf", 
X"7db1", X"7db3", X"7db6", X"7db8", X"7dba", X"7dbd", X"7dbf", X"7dc2", 
X"7dc4", X"7dc6", X"7dc9", X"7dcb", X"7dcd", X"7dcf", X"7dd2", X"7dd4", 
X"7dd6", X"7dd9", X"7ddb", X"7ddd", X"7de0", X"7de2", X"7de4", X"7de6", 
X"7de9", X"7deb", X"7ded", X"7def", X"7df2", X"7df4", X"7df6", X"7df8", 
X"7dfb", X"7dfd", X"7dff", X"7e01", X"7e03", X"7e06", X"7e08", X"7e0a", 
X"7e0c", X"7e0e", X"7e11", X"7e13", X"7e15", X"7e17", X"7e19", X"7e1b", 
X"7e1e", X"7e20", X"7e22", X"7e24", X"7e26", X"7e28", X"7e2a", X"7e2d", 
X"7e2f", X"7e31", X"7e33", X"7e35", X"7e37", X"7e39", X"7e3b", X"7e3d", 
X"7e3f", X"7e41", X"7e43", X"7e46", X"7e48", X"7e4a", X"7e4c", X"7e4e", 
X"7e50", X"7e52", X"7e54", X"7e56", X"7e58", X"7e5a", X"7e5c", X"7e5e", 
X"7e60", X"7e62", X"7e64", X"7e66", X"7e68", X"7e6a", X"7e6c", X"7e6e", 
X"7e70", X"7e72", X"7e74", X"7e76", X"7e78", X"7e79", X"7e7b", X"7e7d", 
X"7e7f", X"7e81", X"7e83", X"7e85", X"7e87", X"7e89", X"7e8b", X"7e8d", 
X"7e8e", X"7e90", X"7e92", X"7e94", X"7e96", X"7e98", X"7e9a", X"7e9b", 
X"7e9d", X"7e9f", X"7ea1", X"7ea3", X"7ea5", X"7ea6", X"7ea8", X"7eaa", 
X"7eac", X"7eae", X"7eb0", X"7eb1", X"7eb3", X"7eb5", X"7eb7", X"7eb8", 
X"7eba", X"7ebc", X"7ebe", X"7ec0", X"7ec1", X"7ec3", X"7ec5", X"7ec6", 
X"7ec8", X"7eca", X"7ecc", X"7ecd", X"7ecf", X"7ed1", X"7ed3", X"7ed4", 
X"7ed6", X"7ed8", X"7ed9", X"7edb", X"7edd", X"7ede", X"7ee0", X"7ee2", 
X"7ee3", X"7ee5", X"7ee7", X"7ee8", X"7eea", X"7eeb", X"7eed", X"7eef", 
X"7ef0", X"7ef2", X"7ef4", X"7ef5", X"7ef7", X"7ef8", X"7efa", X"7efc", 
X"7efd", X"7eff", X"7f00", X"7f02", X"7f03", X"7f05", X"7f06", X"7f08", 
X"7f0a", X"7f0b", X"7f0d", X"7f0e", X"7f10", X"7f11", X"7f13", X"7f14", 
X"7f16", X"7f17", X"7f19", X"7f1a", X"7f1c", X"7f1d", X"7f1f", X"7f20", 
X"7f22", X"7f23", X"7f24", X"7f26", X"7f27", X"7f29", X"7f2a", X"7f2c", 
X"7f2d", X"7f2f", X"7f30", X"7f31", X"7f33", X"7f34", X"7f36", X"7f37", 
X"7f38", X"7f3a", X"7f3b", X"7f3c", X"7f3e", X"7f3f", X"7f41", X"7f42", 
X"7f43", X"7f45", X"7f46", X"7f47", X"7f49", X"7f4a", X"7f4b", X"7f4d", 
X"7f4e", X"7f4f", X"7f50", X"7f52", X"7f53", X"7f54", X"7f56", X"7f57", 
X"7f58", X"7f59", X"7f5b", X"7f5c", X"7f5d", X"7f5e", X"7f60", X"7f61", 
X"7f62", X"7f63", X"7f65", X"7f66", X"7f67", X"7f68", X"7f6a", X"7f6b", 
X"7f6c", X"7f6d", X"7f6e", X"7f6f", X"7f71", X"7f72", X"7f73", X"7f74", 
X"7f75", X"7f76", X"7f78", X"7f79", X"7f7a", X"7f7b", X"7f7c", X"7f7d", 
X"7f7e", X"7f80", X"7f81", X"7f82", X"7f83", X"7f84", X"7f85", X"7f86", 
X"7f87", X"7f88", X"7f89", X"7f8a", X"7f8b", X"7f8d", X"7f8e", X"7f8f", 
X"7f90", X"7f91", X"7f92", X"7f93", X"7f94", X"7f95", X"7f96", X"7f97", 
X"7f98", X"7f99", X"7f9a", X"7f9b", X"7f9c", X"7f9d", X"7f9e", X"7f9f", 
X"7fa0", X"7fa1", X"7fa2", X"7fa3", X"7fa3", X"7fa4", X"7fa5", X"7fa6", 
X"7fa7", X"7fa8", X"7fa9", X"7faa", X"7fab", X"7fac", X"7fad", X"7fae", 
X"7fae", X"7faf", X"7fb0", X"7fb1", X"7fb2", X"7fb3", X"7fb4", X"7fb5", 
X"7fb5", X"7fb6", X"7fb7", X"7fb8", X"7fb9", X"7fba", X"7fba", X"7fbb", 
X"7fbc", X"7fbd", X"7fbe", X"7fbe", X"7fbf", X"7fc0", X"7fc1", X"7fc2", 
X"7fc2", X"7fc3", X"7fc4", X"7fc5", X"7fc5", X"7fc6", X"7fc7", X"7fc8", 
X"7fc8", X"7fc9", X"7fca", X"7fcb", X"7fcb", X"7fcc", X"7fcd", X"7fcd", 
X"7fce", X"7fcf", X"7fcf", X"7fd0", X"7fd1", X"7fd1", X"7fd2", X"7fd3", 
X"7fd3", X"7fd4", X"7fd5", X"7fd5", X"7fd6", X"7fd7", X"7fd7", X"7fd8", 
X"7fd9", X"7fd9", X"7fda", X"7fda", X"7fdb", X"7fdc", X"7fdc", X"7fdd", 
X"7fdd", X"7fde", X"7fde", X"7fdf", X"7fe0", X"7fe0", X"7fe1", X"7fe1", 
X"7fe2", X"7fe2", X"7fe3", X"7fe3", X"7fe4", X"7fe4", X"7fe5", X"7fe5", 
X"7fe6", X"7fe6", X"7fe7", X"7fe7", X"7fe8", X"7fe8", X"7fe9", X"7fe9", 
X"7fea", X"7fea", X"7feb", X"7feb", X"7fec", X"7fec", X"7fec", X"7fed", 
X"7fed", X"7fee", X"7fee", X"7fef", X"7fef", X"7fef", X"7ff0", X"7ff0", 
X"7ff1", X"7ff1", X"7ff1", X"7ff2", X"7ff2", X"7ff2", X"7ff3", X"7ff3", 
X"7ff4", X"7ff4", X"7ff4", X"7ff5", X"7ff5", X"7ff5", X"7ff6", X"7ff6", 
X"7ff6", X"7ff6", X"7ff7", X"7ff7", X"7ff7", X"7ff8", X"7ff8", X"7ff8", 
X"7ff8", X"7ff9", X"7ff9", X"7ff9", X"7ff9", X"7ffa", X"7ffa", X"7ffa", 
X"7ffa", X"7ffb", X"7ffb", X"7ffb", X"7ffb", X"7ffc", X"7ffc", X"7ffc", 
X"7ffc", X"7ffc", X"7ffd", X"7ffd", X"7ffd", X"7ffd", X"7ffd", X"7ffd", 
X"7ffe", X"7ffe", X"7ffe", X"7ffe", X"7ffe", X"7ffe", X"7ffe", X"7ffe", 
X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", 
X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", 
X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", 
X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", 
X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", 
X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", X"7fff", 
X"7fff", X"7ffe", X"7ffe", X"7ffe", X"7ffe", X"7ffe", X"7ffe", X"7ffe", 
X"7ffe", X"7ffd", X"7ffd", X"7ffd", X"7ffd", X"7ffd", X"7ffd", X"7ffc", 
X"7ffc", X"7ffc", X"7ffc", X"7ffc", X"7ffb", X"7ffb", X"7ffb", X"7ffb", 
X"7ffa", X"7ffa", X"7ffa", X"7ffa", X"7ff9", X"7ff9", X"7ff9", X"7ff9", 
X"7ff8", X"7ff8", X"7ff8", X"7ff8", X"7ff7", X"7ff7", X"7ff7", X"7ff6", 
X"7ff6", X"7ff6", X"7ff6", X"7ff5", X"7ff5", X"7ff5", X"7ff4", X"7ff4", 
X"7ff4", X"7ff3", X"7ff3", X"7ff2", X"7ff2", X"7ff2", X"7ff1", X"7ff1", 
X"7ff1", X"7ff0", X"7ff0", X"7fef", X"7fef", X"7fef", X"7fee", X"7fee", 
X"7fed", X"7fed", X"7fec", X"7fec", X"7fec", X"7feb", X"7feb", X"7fea", 
X"7fea", X"7fe9", X"7fe9", X"7fe8", X"7fe8", X"7fe7", X"7fe7", X"7fe6", 
X"7fe6", X"7fe5", X"7fe5", X"7fe4", X"7fe4", X"7fe3", X"7fe3", X"7fe2", 
X"7fe2", X"7fe1", X"7fe1", X"7fe0", X"7fe0", X"7fdf", X"7fde", X"7fde", 
X"7fdd", X"7fdd", X"7fdc", X"7fdc", X"7fdb", X"7fda", X"7fda", X"7fd9", 
X"7fd9", X"7fd8", X"7fd7", X"7fd7", X"7fd6", X"7fd5", X"7fd5", X"7fd4", 
X"7fd3", X"7fd3", X"7fd2", X"7fd1", X"7fd1", X"7fd0", X"7fcf", X"7fcf", 
X"7fce", X"7fcd", X"7fcd", X"7fcc", X"7fcb", X"7fcb", X"7fca", X"7fc9", 
X"7fc8", X"7fc8", X"7fc7", X"7fc6", X"7fc5", X"7fc5", X"7fc4", X"7fc3", 
X"7fc2", X"7fc2", X"7fc1", X"7fc0", X"7fbf", X"7fbe", X"7fbe", X"7fbd", 
X"7fbc", X"7fbb", X"7fba", X"7fba", X"7fb9", X"7fb8", X"7fb7", X"7fb6", 
X"7fb5", X"7fb5", X"7fb4", X"7fb3", X"7fb2", X"7fb1", X"7fb0", X"7faf", 
X"7fae", X"7fae", X"7fad", X"7fac", X"7fab", X"7faa", X"7fa9", X"7fa8", 
X"7fa7", X"7fa6", X"7fa5", X"7fa4", X"7fa3", X"7fa3", X"7fa2", X"7fa1", 
X"7fa0", X"7f9f", X"7f9e", X"7f9d", X"7f9c", X"7f9b", X"7f9a", X"7f99", 
X"7f98", X"7f97", X"7f96", X"7f95", X"7f94", X"7f93", X"7f92", X"7f91", 
X"7f90", X"7f8f", X"7f8e", X"7f8d", X"7f8b", X"7f8a", X"7f89", X"7f88", 
X"7f87", X"7f86", X"7f85", X"7f84", X"7f83", X"7f82", X"7f81", X"7f80", 
X"7f7e", X"7f7d", X"7f7c", X"7f7b", X"7f7a", X"7f79", X"7f78", X"7f76", 
X"7f75", X"7f74", X"7f73", X"7f72", X"7f71", X"7f6f", X"7f6e", X"7f6d", 
X"7f6c", X"7f6b", X"7f6a", X"7f68", X"7f67", X"7f66", X"7f65", X"7f63", 
X"7f62", X"7f61", X"7f60", X"7f5e", X"7f5d", X"7f5c", X"7f5b", X"7f59", 
X"7f58", X"7f57", X"7f56", X"7f54", X"7f53", X"7f52", X"7f50", X"7f4f", 
X"7f4e", X"7f4d", X"7f4b", X"7f4a", X"7f49", X"7f47", X"7f46", X"7f45", 
X"7f43", X"7f42", X"7f41", X"7f3f", X"7f3e", X"7f3c", X"7f3b", X"7f3a", 
X"7f38", X"7f37", X"7f36", X"7f34", X"7f33", X"7f31", X"7f30", X"7f2f", 
X"7f2d", X"7f2c", X"7f2a", X"7f29", X"7f27", X"7f26", X"7f24", X"7f23", 
X"7f22", X"7f20", X"7f1f", X"7f1d", X"7f1c", X"7f1a", X"7f19", X"7f17", 
X"7f16", X"7f14", X"7f13", X"7f11", X"7f10", X"7f0e", X"7f0d", X"7f0b", 
X"7f0a", X"7f08", X"7f06", X"7f05", X"7f03", X"7f02", X"7f00", X"7eff", 
X"7efd", X"7efc", X"7efa", X"7ef8", X"7ef7", X"7ef5", X"7ef4", X"7ef2", 
X"7ef0", X"7eef", X"7eed", X"7eeb", X"7eea", X"7ee8", X"7ee7", X"7ee5", 
X"7ee3", X"7ee2", X"7ee0", X"7ede", X"7edd", X"7edb", X"7ed9", X"7ed8", 
X"7ed6", X"7ed4", X"7ed3", X"7ed1", X"7ecf", X"7ecd", X"7ecc", X"7eca", 
X"7ec8", X"7ec6", X"7ec5", X"7ec3", X"7ec1", X"7ec0", X"7ebe", X"7ebc", 
X"7eba", X"7eb8", X"7eb7", X"7eb5", X"7eb3", X"7eb1", X"7eb0", X"7eae", 
X"7eac", X"7eaa", X"7ea8", X"7ea6", X"7ea5", X"7ea3", X"7ea1", X"7e9f", 
X"7e9d", X"7e9b", X"7e9a", X"7e98", X"7e96", X"7e94", X"7e92", X"7e90", 
X"7e8e", X"7e8d", X"7e8b", X"7e89", X"7e87", X"7e85", X"7e83", X"7e81", 
X"7e7f", X"7e7d", X"7e7b", X"7e79", X"7e78", X"7e76", X"7e74", X"7e72", 
X"7e70", X"7e6e", X"7e6c", X"7e6a", X"7e68", X"7e66", X"7e64", X"7e62", 
X"7e60", X"7e5e", X"7e5c", X"7e5a", X"7e58", X"7e56", X"7e54", X"7e52", 
X"7e50", X"7e4e", X"7e4c", X"7e4a", X"7e48", X"7e46", X"7e43", X"7e41", 
X"7e3f", X"7e3d", X"7e3b", X"7e39", X"7e37", X"7e35", X"7e33", X"7e31", 
X"7e2f", X"7e2d", X"7e2a", X"7e28", X"7e26", X"7e24", X"7e22", X"7e20", 
X"7e1e", X"7e1b", X"7e19", X"7e17", X"7e15", X"7e13", X"7e11", X"7e0e", 
X"7e0c", X"7e0a", X"7e08", X"7e06", X"7e03", X"7e01", X"7dff", X"7dfd", 
X"7dfb", X"7df8", X"7df6", X"7df4", X"7df2", X"7def", X"7ded", X"7deb", 
X"7de9", X"7de6", X"7de4", X"7de2", X"7de0", X"7ddd", X"7ddb", X"7dd9", 
X"7dd6", X"7dd4", X"7dd2", X"7dcf", X"7dcd", X"7dcb", X"7dc9", X"7dc6", 
X"7dc4", X"7dc2", X"7dbf", X"7dbd", X"7dba", X"7db8", X"7db6", X"7db3", 
X"7db1", X"7daf", X"7dac", X"7daa", X"7da7", X"7da5", X"7da3", X"7da0", 
X"7d9e", X"7d9b", X"7d99", X"7d97", X"7d94", X"7d92", X"7d8f", X"7d8d", 
X"7d8a", X"7d88", X"7d85", X"7d83", X"7d81", X"7d7e", X"7d7c", X"7d79", 
X"7d77", X"7d74", X"7d72", X"7d6f", X"7d6d", X"7d6a", X"7d68", X"7d65", 
X"7d63", X"7d60", X"7d5d", X"7d5b", X"7d58", X"7d56", X"7d53", X"7d51", 
X"7d4e", X"7d4c", X"7d49", X"7d46", X"7d44", X"7d41", X"7d3f", X"7d3c", 
X"7d3a", X"7d37", X"7d34", X"7d32", X"7d2f", X"7d2c", X"7d2a", X"7d27", 
X"7d25", X"7d22", X"7d1f", X"7d1d", X"7d1a", X"7d17", X"7d15", X"7d12", 
X"7d0f", X"7d0d", X"7d0a", X"7d07", X"7d05", X"7d02", X"7cff", X"7cfc", 
X"7cfa", X"7cf7", X"7cf4", X"7cf2", X"7cef", X"7cec", X"7ce9", X"7ce7", 
X"7ce4", X"7ce1", X"7cde", X"7cdc", X"7cd9", X"7cd6", X"7cd3", X"7cd0", 
X"7cce", X"7ccb", X"7cc8", X"7cc5", X"7cc2", X"7cc0", X"7cbd", X"7cba", 
X"7cb7", X"7cb4", X"7cb1", X"7caf", X"7cac", X"7ca9", X"7ca6", X"7ca3", 
X"7ca0", X"7c9e", X"7c9b", X"7c98", X"7c95", X"7c92", X"7c8f", X"7c8c", 
X"7c89", X"7c86", X"7c83", X"7c81", X"7c7e", X"7c7b", X"7c78", X"7c75", 
X"7c72", X"7c6f", X"7c6c", X"7c69", X"7c66", X"7c63", X"7c60", X"7c5d", 
X"7c5a", X"7c57", X"7c54", X"7c51", X"7c4e", X"7c4b", X"7c48", X"7c45", 
X"7c42", X"7c3f", X"7c3c", X"7c39", X"7c36", X"7c33", X"7c30", X"7c2d", 
X"7c2a", X"7c27", X"7c24", X"7c21", X"7c1e", X"7c1b", X"7c18", X"7c14", 
X"7c11", X"7c0e", X"7c0b", X"7c08", X"7c05", X"7c02", X"7bff", X"7bfc", 
X"7bf9", X"7bf5", X"7bf2", X"7bef", X"7bec", X"7be9", X"7be6", X"7be3", 
X"7bdf", X"7bdc", X"7bd9", X"7bd6", X"7bd3", X"7bcf", X"7bcc", X"7bc9", 
X"7bc6", X"7bc3", X"7bbf", X"7bbc", X"7bb9", X"7bb6", X"7bb3", X"7baf", 
X"7bac", X"7ba9", X"7ba6", X"7ba2", X"7b9f", X"7b9c", X"7b99", X"7b95", 
X"7b92", X"7b8f", X"7b8b", X"7b88", X"7b85", X"7b82", X"7b7e", X"7b7b", 
X"7b78", X"7b74", X"7b71", X"7b6e", X"7b6a", X"7b67", X"7b64", X"7b60", 
X"7b5d", X"7b5a", X"7b56", X"7b53", X"7b50", X"7b4c", X"7b49", X"7b45", 
X"7b42", X"7b3f", X"7b3b", X"7b38", X"7b34", X"7b31", X"7b2e", X"7b2a", 
X"7b27", X"7b23", X"7b20", X"7b1c", X"7b19", X"7b16", X"7b12", X"7b0f", 
X"7b0b", X"7b08", X"7b04", X"7b01", X"7afd", X"7afa", X"7af6", X"7af3", 
X"7aef", X"7aec", X"7ae8", X"7ae5", X"7ae1", X"7ade", X"7ada", X"7ad7", 
X"7ad3", X"7ad0", X"7acc", X"7ac9", X"7ac5", X"7ac1", X"7abe", X"7aba", 
X"7ab7", X"7ab3", X"7ab0", X"7aac", X"7aa8", X"7aa5", X"7aa1", X"7a9e", 
X"7a9a", X"7a96", X"7a93", X"7a8f", X"7a8c", X"7a88", X"7a84", X"7a81", 
X"7a7d", X"7a79", X"7a76", X"7a72", X"7a6e", X"7a6b", X"7a67", X"7a63", 
X"7a60", X"7a5c", X"7a58", X"7a55", X"7a51", X"7a4d", X"7a49", X"7a46", 
X"7a42", X"7a3e", X"7a3b", X"7a37", X"7a33", X"7a2f", X"7a2c", X"7a28", 
X"7a24", X"7a20", X"7a1d", X"7a19", X"7a15", X"7a11", X"7a0e", X"7a0a", 
X"7a06", X"7a02", X"79fe", X"79fb", X"79f7", X"79f3", X"79ef", X"79eb", 
X"79e7", X"79e4", X"79e0", X"79dc", X"79d8", X"79d4", X"79d0", X"79cc", 
X"79c9", X"79c5", X"79c1", X"79bd", X"79b9", X"79b5", X"79b1", X"79ad", 
X"79aa", X"79a6", X"79a2", X"799e", X"799a", X"7996", X"7992", X"798e", 
X"798a", X"7986", X"7982", X"797e", X"797a", X"7976", X"7972", X"796e", 
X"796a", X"7966", X"7962", X"795f", X"795b", X"7957", X"7953", X"794e", 
X"794a", X"7946", X"7942", X"793e", X"793a", X"7936", X"7932", X"792e", 
X"792a", X"7926", X"7922", X"791e", X"791a", X"7916", X"7912", X"790e", 
X"790a", X"7906", X"7901", X"78fd", X"78f9", X"78f5", X"78f1", X"78ed", 
X"78e9", X"78e5", X"78e1", X"78dc", X"78d8", X"78d4", X"78d0", X"78cc", 
X"78c8", X"78c4", X"78bf", X"78bb", X"78b7", X"78b3", X"78af", X"78aa", 
X"78a6", X"78a2", X"789e", X"789a", X"7895", X"7891", X"788d", X"7889", 
X"7885", X"7880", X"787c", X"7878", X"7874", X"786f", X"786b", X"7867", 
X"7863", X"785e", X"785a", X"7856", X"7851", X"784d", X"7849", X"7845", 
X"7840", X"783c", X"7838", X"7833", X"782f", X"782b", X"7826", X"7822", 
X"781e", X"7819", X"7815", X"7811", X"780c", X"7808", X"7803", X"77ff", 
X"77fb", X"77f6", X"77f2", X"77ee", X"77e9", X"77e5", X"77e0", X"77dc", 
X"77d8", X"77d3", X"77cf", X"77ca", X"77c6", X"77c1", X"77bd", X"77b9", 
X"77b4", X"77b0", X"77ab", X"77a7", X"77a2", X"779e", X"7799", X"7795", 
X"7790", X"778c", X"7787", X"7783", X"777e", X"777a", X"7775", X"7771", 
X"776c", X"7768", X"7763", X"775f", X"775a", X"7756", X"7751", X"774d", 
X"7748", X"7743", X"773f", X"773a", X"7736", X"7731", X"772d", X"7728", 
X"7723", X"771f", X"771a", X"7716", X"7711", X"770c", X"7708", X"7703", 
X"76fe", X"76fa", X"76f5", X"76f1", X"76ec", X"76e7", X"76e3", X"76de", 
X"76d9", X"76d5", X"76d0", X"76cb", X"76c7", X"76c2", X"76bd", X"76b9", 
X"76b4", X"76af", X"76aa", X"76a6", X"76a1", X"769c", X"7698", X"7693", 
X"768e", X"7689", X"7685", X"7680", X"767b", X"7676", X"7672", X"766d", 
X"7668", X"7663", X"765e", X"765a", X"7655", X"7650", X"764b", X"7646", 
X"7642", X"763d", X"7638", X"7633", X"762e", X"762a", X"7625", X"7620", 
X"761b", X"7616", X"7611", X"760d", X"7608", X"7603", X"75fe", X"75f9", 
X"75f4", X"75ef", X"75ea", X"75e6", X"75e1", X"75dc", X"75d7", X"75d2", 
X"75cd", X"75c8", X"75c3", X"75be", X"75b9", X"75b4", X"75af", X"75aa", 
X"75a6", X"75a1", X"759c", X"7597", X"7592", X"758d", X"7588", X"7583", 
X"757e", X"7579", X"7574", X"756f", X"756a", X"7565", X"7560", X"755b", 
X"7556", X"7551", X"754c", X"7547", X"7542", X"753d", X"7538", X"7532", 
X"752d", X"7528", X"7523", X"751e", X"7519", X"7514", X"750f", X"750a", 
X"7505", X"7500", X"74fb", X"74f6", X"74f0", X"74eb", X"74e6", X"74e1", 
X"74dc", X"74d7", X"74d2", X"74cd", X"74c7", X"74c2", X"74bd", X"74b8", 
X"74b3", X"74ae", X"74a8", X"74a3", X"749e", X"7499", X"7494", X"748f", 
X"7489", X"7484", X"747f", X"747a", X"7475", X"746f", X"746a", X"7465", 
X"7460", X"745a", X"7455", X"7450", X"744b", X"7445", X"7440", X"743b", 
X"7436", X"7430", X"742b", X"7426", X"7421", X"741b", X"7416", X"7411", 
X"740b", X"7406", X"7401", X"73fb", X"73f6", X"73f1", X"73eb", X"73e6", 
X"73e1", X"73db", X"73d6", X"73d1", X"73cb", X"73c6", X"73c1", X"73bb", 
X"73b6", X"73b1", X"73ab", X"73a6", X"73a0", X"739b", X"7396", X"7390", 
X"738b", X"7385", X"7380", X"737b", X"7375", X"7370", X"736a", X"7365", 
X"735f", X"735a", X"7355", X"734f", X"734a", X"7344", X"733f", X"7339", 
X"7334", X"732e", X"7329", X"7323", X"731e", X"7318", X"7313", X"730d", 
X"7308", X"7302", X"72fd", X"72f7", X"72f2", X"72ec", X"72e7", X"72e1", 
X"72dc", X"72d6", X"72d0", X"72cb", X"72c5", X"72c0", X"72ba", X"72b5", 
X"72af", X"72a9", X"72a4", X"729e", X"7299", X"7293", X"728d", X"7288", 
X"7282", X"727d", X"7277", X"7271", X"726c", X"7266", X"7260", X"725b", 
X"7255", X"7250", X"724a", X"7244", X"723f", X"7239", X"7233", X"722e", 
X"7228", X"7222", X"721c", X"7217", X"7211", X"720b", X"7206", X"7200", 
X"71fa", X"71f5", X"71ef", X"71e9", X"71e3", X"71de", X"71d8", X"71d2", 
X"71cc", X"71c7", X"71c1", X"71bb", X"71b5", X"71b0", X"71aa", X"71a4", 
X"719e", X"7198", X"7193", X"718d", X"7187", X"7181", X"717b", X"7176", 
X"7170", X"716a", X"7164", X"715e", X"7158", X"7153", X"714d", X"7147", 
X"7141", X"713b", X"7135", X"712f", X"712a", X"7124", X"711e", X"7118", 
X"7112", X"710c", X"7106", X"7100", X"70fa", X"70f5", X"70ef", X"70e9", 
X"70e3", X"70dd", X"70d7", X"70d1", X"70cb", X"70c5", X"70bf", X"70b9", 
X"70b3", X"70ad", X"70a7", X"70a1", X"709b", X"7095", X"708f", X"7089", 
X"7083", X"707d", X"7077", X"7071", X"706b", X"7065", X"705f", X"7059", 
X"7053", X"704d", X"7047", X"7041", X"703b", X"7035", X"702f", X"7029", 
X"7023", X"701d", X"7017", X"7011", X"700b", X"7005", X"6fff", X"6ff9", 
X"6ff2", X"6fec", X"6fe6", X"6fe0", X"6fda", X"6fd4", X"6fce", X"6fc8", 
X"6fc2", X"6fbb", X"6fb5", X"6faf", X"6fa9", X"6fa3", X"6f9d", X"6f97", 
X"6f90", X"6f8a", X"6f84", X"6f7e", X"6f78", X"6f72", X"6f6b", X"6f65", 
X"6f5f", X"6f59", X"6f53", X"6f4c", X"6f46", X"6f40", X"6f3a", X"6f34", 
X"6f2d", X"6f27", X"6f21", X"6f1b", X"6f14", X"6f0e", X"6f08", X"6f02", 
X"6efb", X"6ef5", X"6eef", X"6ee9", X"6ee2", X"6edc", X"6ed6", X"6ecf", 
X"6ec9", X"6ec3", X"6ebd", X"6eb6", X"6eb0", X"6eaa", X"6ea3", X"6e9d", 
X"6e97", X"6e90", X"6e8a", X"6e84", X"6e7d", X"6e77", X"6e71", X"6e6a", 
X"6e64", X"6e5e", X"6e57", X"6e51", X"6e4a", X"6e44", X"6e3e", X"6e37", 
X"6e31", X"6e2a", X"6e24", X"6e1e", X"6e17", X"6e11", X"6e0a", X"6e04", 
X"6dfe", X"6df7", X"6df1", X"6dea", X"6de4", X"6ddd", X"6dd7", X"6dd1", 
X"6dca", X"6dc4", X"6dbd", X"6db7", X"6db0", X"6daa", X"6da3", X"6d9d", 
X"6d96", X"6d90", X"6d89", X"6d83", X"6d7c", X"6d76", X"6d6f", X"6d69", 
X"6d62", X"6d5c", X"6d55", X"6d4f", X"6d48", X"6d41", X"6d3b", X"6d34", 
X"6d2e", X"6d27", X"6d21", X"6d1a", X"6d14", X"6d0d", X"6d06", X"6d00", 
X"6cf9", X"6cf3", X"6cec", X"6ce5", X"6cdf", X"6cd8", X"6cd2", X"6ccb", 
X"6cc4", X"6cbe", X"6cb7", X"6cb0", X"6caa", X"6ca3", X"6c9d", X"6c96", 
X"6c8f", X"6c89", X"6c82", X"6c7b", X"6c75", X"6c6e", X"6c67", X"6c61", 
X"6c5a", X"6c53", X"6c4c", X"6c46", X"6c3f", X"6c38", X"6c32", X"6c2b", 
X"6c24", X"6c1d", X"6c17", X"6c10", X"6c09", X"6c02", X"6bfc", X"6bf5", 
X"6bee", X"6be7", X"6be1", X"6bda", X"6bd3", X"6bcc", X"6bc6", X"6bbf", 
X"6bb8", X"6bb1", X"6baa", X"6ba4", X"6b9d", X"6b96", X"6b8f", X"6b88", 
X"6b82", X"6b7b", X"6b74", X"6b6d", X"6b66", X"6b5f", X"6b59", X"6b52", 
X"6b4b", X"6b44", X"6b3d", X"6b36", X"6b30", X"6b29", X"6b22", X"6b1b", 
X"6b14", X"6b0d", X"6b06", X"6aff", X"6af8", X"6af2", X"6aeb", X"6ae4", 
X"6add", X"6ad6", X"6acf", X"6ac8", X"6ac1", X"6aba", X"6ab3", X"6aac", 
X"6aa5", X"6a9e", X"6a97", X"6a90", X"6a89", X"6a83", X"6a7c", X"6a75", 
X"6a6e", X"6a67", X"6a60", X"6a59", X"6a52", X"6a4b", X"6a44", X"6a3d", 
X"6a36", X"6a2f", X"6a28", X"6a21", X"6a1a", X"6a12", X"6a0b", X"6a04", 
X"69fd", X"69f6", X"69ef", X"69e8", X"69e1", X"69da", X"69d3", X"69cc", 
X"69c5", X"69be", X"69b7", X"69b0", X"69a9", X"69a1", X"699a", X"6993", 
X"698c", X"6985", X"697e", X"6977", X"6970", X"6969", X"6961", X"695a", 
X"6953", X"694c", X"6945", X"693e", X"6937", X"692f", X"6928", X"6921", 
X"691a", X"6913", X"690c", X"6904", X"68fd", X"68f6", X"68ef", X"68e8", 
X"68e0", X"68d9", X"68d2", X"68cb", X"68c4", X"68bc", X"68b5", X"68ae", 
X"68a7", X"689f", X"6898", X"6891", X"688a", X"6882", X"687b", X"6874", 
X"686d", X"6865", X"685e", X"6857", X"6850", X"6848", X"6841", X"683a", 
X"6832", X"682b", X"6824", X"681c", X"6815", X"680e", X"6806", X"67ff", 
X"67f8", X"67f0", X"67e9", X"67e2", X"67da", X"67d3", X"67cc", X"67c4", 
X"67bd", X"67b6", X"67ae", X"67a7", X"67a0", X"6798", X"6791", X"6789", 
X"6782", X"677b", X"6773", X"676c", X"6764", X"675d", X"6756", X"674e", 
X"6747", X"673f", X"6738", X"6730", X"6729", X"6722", X"671a", X"6713", 
X"670b", X"6704", X"66fc", X"66f5", X"66ed", X"66e6", X"66de", X"66d7", 
X"66d0", X"66c8", X"66c1", X"66b9", X"66b2", X"66aa", X"66a3", X"669b", 
X"6693", X"668c", X"6684", X"667d", X"6675", X"666e", X"6666", X"665f", 
X"6657", X"6650", X"6648", X"6641", X"6639", X"6631", X"662a", X"6622", 
X"661b", X"6613", X"660c", X"6604", X"65fc", X"65f5", X"65ed", X"65e6", 
X"65de", X"65d6", X"65cf", X"65c7", X"65c0", X"65b8", X"65b0", X"65a9", 
X"65a1", X"6599", X"6592", X"658a", X"6582", X"657b", X"6573", X"656b", 
X"6564", X"655c", X"6554", X"654d", X"6545", X"653d", X"6536", X"652e", 
X"6526", X"651f", X"6517", X"650f", X"6507", X"6500", X"64f8", X"64f0", 
X"64e9", X"64e1", X"64d9", X"64d1", X"64ca", X"64c2", X"64ba", X"64b2", 
X"64ab", X"64a3", X"649b", X"6493", X"648b", X"6484", X"647c", X"6474", 
X"646c", X"6465", X"645d", X"6455", X"644d", X"6445", X"643e", X"6436", 
X"642e", X"6426", X"641e", X"6416", X"640f", X"6407", X"63ff", X"63f7", 
X"63ef", X"63e7", X"63df", X"63d8", X"63d0", X"63c8", X"63c0", X"63b8", 
X"63b0", X"63a8", X"63a0", X"6399", X"6391", X"6389", X"6381", X"6379", 
X"6371", X"6369", X"6361", X"6359", X"6351", X"6349", X"6342", X"633a", 
X"6332", X"632a", X"6322", X"631a", X"6312", X"630a", X"6302", X"62fa", 
X"62f2", X"62ea", X"62e2", X"62da", X"62d2", X"62ca", X"62c2", X"62ba", 
X"62b2", X"62aa", X"62a2", X"629a", X"6292", X"628a", X"6282", X"627a", 
X"6272", X"626a", X"6262", X"625a", X"6252", X"624a", X"6242", X"623a", 
X"6232", X"622a", X"6221", X"6219", X"6211", X"6209", X"6201", X"61f9", 
X"61f1", X"61e9", X"61e1", X"61d9", X"61d1", X"61c9", X"61c0", X"61b8", 
X"61b0", X"61a8", X"61a0", X"6198", X"6190", X"6188", X"617f", X"6177", 
X"616f", X"6167", X"615f", X"6157", X"614e", X"6146", X"613e", X"6136", 
X"612e", X"6126", X"611d", X"6115", X"610d", X"6105", X"60fd", X"60f4", 
X"60ec", X"60e4", X"60dc", X"60d4", X"60cb", X"60c3", X"60bb", X"60b3", 
X"60aa", X"60a2", X"609a", X"6092", X"6089", X"6081", X"6079", X"6071", 
X"6068", X"6060", X"6058", X"6050", X"6047", X"603f", X"6037", X"602e", 
X"6026", X"601e", X"6016", X"600d", X"6005", X"5ffd", X"5ff4", X"5fec", 
X"5fe4", X"5fdb", X"5fd3", X"5fcb", X"5fc2", X"5fba", X"5fb2", X"5fa9", 
X"5fa1", X"5f99", X"5f90", X"5f88", X"5f80", X"5f77", X"5f6f", X"5f66", 
X"5f5e", X"5f56", X"5f4d", X"5f45", X"5f3c", X"5f34", X"5f2c", X"5f23", 
X"5f1b", X"5f12", X"5f0a", X"5f02", X"5ef9", X"5ef1", X"5ee8", X"5ee0", 
X"5ed7", X"5ecf", X"5ec7", X"5ebe", X"5eb6", X"5ead", X"5ea5", X"5e9c", 
X"5e94", X"5e8b", X"5e83", X"5e7a", X"5e72", X"5e69", X"5e61", X"5e58", 
X"5e50", X"5e48", X"5e3f", X"5e37", X"5e2e", X"5e25", X"5e1d", X"5e14", 
X"5e0c", X"5e03", X"5dfb", X"5df2", X"5dea", X"5de1", X"5dd9", X"5dd0", 
X"5dc8", X"5dbf", X"5db7", X"5dae", X"5da5", X"5d9d", X"5d94", X"5d8c", 
X"5d83", X"5d7a", X"5d72", X"5d69", X"5d61", X"5d58", X"5d50", X"5d47", 
X"5d3e", X"5d36", X"5d2d", X"5d24", X"5d1c", X"5d13", X"5d0b", X"5d02", 
X"5cf9", X"5cf1", X"5ce8", X"5cdf", X"5cd7", X"5cce", X"5cc5", X"5cbd", 
X"5cb4", X"5cab", X"5ca3", X"5c9a", X"5c91", X"5c89", X"5c80", X"5c77", 
X"5c6f", X"5c66", X"5c5d", X"5c55", X"5c4c", X"5c43", X"5c3a", X"5c32", 
X"5c29", X"5c20", X"5c18", X"5c0f", X"5c06", X"5bfd", X"5bf5", X"5bec", 
X"5be3", X"5bda", X"5bd2", X"5bc9", X"5bc0", X"5bb7", X"5baf", X"5ba6", 
X"5b9d", X"5b94", X"5b8c", X"5b83", X"5b7a", X"5b71", X"5b68", X"5b60", 
X"5b57", X"5b4e", X"5b45", X"5b3c", X"5b34", X"5b2b", X"5b22", X"5b19", 
X"5b10", X"5b07", X"5aff", X"5af6", X"5aed", X"5ae4", X"5adb", X"5ad2", 
X"5ac9", X"5ac1", X"5ab8", X"5aaf", X"5aa6", X"5a9d", X"5a94", X"5a8b", 
X"5a82", X"5a7a", X"5a71", X"5a68", X"5a5f", X"5a56", X"5a4d", X"5a44", 
X"5a3b", X"5a32", X"5a29", X"5a21", X"5a18", X"5a0f", X"5a06", X"59fd", 
X"59f4", X"59eb", X"59e2", X"59d9", X"59d0", X"59c7", X"59be", X"59b5", 
X"59ac", X"59a3", X"599a", X"5991", X"5988", X"597f", X"5976", X"596d", 
X"5964", X"595b", X"5952", X"5949", X"5940", X"5937", X"592e", X"5925", 
X"591c", X"5913", X"590a", X"5901", X"58f8", X"58ef", X"58e6", X"58dd", 
X"58d4", X"58cb", X"58c2", X"58b9", X"58b0", X"58a7", X"589e", X"5895", 
X"588c", X"5882", X"5879", X"5870", X"5867", X"585e", X"5855", X"584c", 
X"5843", X"583a", X"5831", X"5828", X"581e", X"5815", X"580c", X"5803", 
X"57fa", X"57f1", X"57e8", X"57df", X"57d5", X"57cc", X"57c3", X"57ba", 
X"57b1", X"57a8", X"579f", X"5795", X"578c", X"5783", X"577a", X"5771", 
X"5767", X"575e", X"5755", X"574c", X"5743", X"573a", X"5730", X"5727", 
X"571e", X"5715", X"570c", X"5702", X"56f9", X"56f0", X"56e7", X"56dd", 
X"56d4", X"56cb", X"56c2", X"56b8", X"56af", X"56a6", X"569d", X"5693", 
X"568a", X"5681", X"5678", X"566e", X"5665", X"565c", X"5653", X"5649", 
X"5640", X"5637", X"562d", X"5624", X"561b", X"5612", X"5608", X"55ff", 
X"55f6", X"55ec", X"55e3", X"55da", X"55d0", X"55c7", X"55be", X"55b4", 
X"55ab", X"55a2", X"5598", X"558f", X"5586", X"557c", X"5573", X"556a", 
X"5560", X"5557", X"554e", X"5544", X"553b", X"5531", X"5528", X"551f", 
X"5515", X"550c", X"5502", X"54f9", X"54f0", X"54e6", X"54dd", X"54d3", 
X"54ca", X"54c1", X"54b7", X"54ae", X"54a4", X"549b", X"5491", X"5488", 
X"547f", X"5475", X"546c", X"5462", X"5459", X"544f", X"5446", X"543c", 
X"5433", X"542a", X"5420", X"5417", X"540d", X"5404", X"53fa", X"53f1", 
X"53e7", X"53de", X"53d4", X"53cb", X"53c1", X"53b8", X"53ae", X"53a5", 
X"539b", X"5392", X"5388", X"537f", X"5375", X"536c", X"5362", X"5358", 
X"534f", X"5345", X"533c", X"5332", X"5329", X"531f", X"5316", X"530c", 
X"5303", X"52f9", X"52ef", X"52e6", X"52dc", X"52d3", X"52c9", X"52bf", 
X"52b6", X"52ac", X"52a3", X"5299", X"5290", X"5286", X"527c", X"5273", 
X"5269", X"525f", X"5256", X"524c", X"5243", X"5239", X"522f", X"5226", 
X"521c", X"5212", X"5209", X"51ff", X"51f5", X"51ec", X"51e2", X"51d8", 
X"51cf", X"51c5", X"51bb", X"51b2", X"51a8", X"519e", X"5195", X"518b", 
X"5181", X"5178", X"516e", X"5164", X"515b", X"5151", X"5147", X"513e", 
X"5134", X"512a", X"5120", X"5117", X"510d", X"5103", X"50f9", X"50f0", 
X"50e6", X"50dc", X"50d3", X"50c9", X"50bf", X"50b5", X"50ac", X"50a2", 
X"5098", X"508e", X"5084", X"507b", X"5071", X"5067", X"505d", X"5054", 
X"504a", X"5040", X"5036", X"502c", X"5023", X"5019", X"500f", X"5005", 
X"4ffb", X"4ff2", X"4fe8", X"4fde", X"4fd4", X"4fca", X"4fc0", X"4fb7", 
X"4fad", X"4fa3", X"4f99", X"4f8f", X"4f85", X"4f7c", X"4f72", X"4f68", 
X"4f5e", X"4f54", X"4f4a", X"4f40", X"4f37", X"4f2d", X"4f23", X"4f19", 
X"4f0f", X"4f05", X"4efb", X"4ef1", X"4ee8", X"4ede", X"4ed4", X"4eca", 
X"4ec0", X"4eb6", X"4eac", X"4ea2", X"4e98", X"4e8e", X"4e84", X"4e7a", 
X"4e71", X"4e67", X"4e5d", X"4e53", X"4e49", X"4e3f", X"4e35", X"4e2b", 
X"4e21", X"4e17", X"4e0d", X"4e03", X"4df9", X"4def", X"4de5", X"4ddb", 
X"4dd1", X"4dc7", X"4dbd", X"4db3", X"4da9", X"4d9f", X"4d95", X"4d8b", 
X"4d81", X"4d77", X"4d6d", X"4d63", X"4d59", X"4d4f", X"4d45", X"4d3b", 
X"4d31", X"4d27", X"4d1d", X"4d13", X"4d09", X"4cff", X"4cf5", X"4ceb", 
X"4ce1", X"4cd7", X"4ccd", X"4cc3", X"4cb9", X"4caf", X"4ca5", X"4c9b", 
X"4c91", X"4c86", X"4c7c", X"4c72", X"4c68", X"4c5e", X"4c54", X"4c4a", 
X"4c40", X"4c36", X"4c2c", X"4c22", X"4c17", X"4c0d", X"4c03", X"4bf9", 
X"4bef", X"4be5", X"4bdb", X"4bd1", X"4bc7", X"4bbc", X"4bb2", X"4ba8", 
X"4b9e", X"4b94", X"4b8a", X"4b80", X"4b75", X"4b6b", X"4b61", X"4b57", 
X"4b4d", X"4b43", X"4b38", X"4b2e", X"4b24", X"4b1a", X"4b10", X"4b06", 
X"4afb", X"4af1", X"4ae7", X"4add", X"4ad3", X"4ac8", X"4abe", X"4ab4", 
X"4aaa", X"4aa0", X"4a95", X"4a8b", X"4a81", X"4a77", X"4a6d", X"4a62", 
X"4a58", X"4a4e", X"4a44", X"4a39", X"4a2f", X"4a25", X"4a1b", X"4a10", 
X"4a06", X"49fc", X"49f2", X"49e7", X"49dd", X"49d3", X"49c9", X"49be", 
X"49b4", X"49aa", X"49a0", X"4995", X"498b", X"4981", X"4976", X"496c", 
X"4962", X"4958", X"494d", X"4943", X"4939", X"492e", X"4924", X"491a", 
X"490f", X"4905", X"48fb", X"48f0", X"48e6", X"48dc", X"48d1", X"48c7", 
X"48bd", X"48b2", X"48a8", X"489e", X"4893", X"4889", X"487f", X"4874", 
X"486a", X"4860", X"4855", X"484b", X"4840", X"4836", X"482c", X"4821", 
X"4817", X"480d", X"4802", X"47f8", X"47ed", X"47e3", X"47d9", X"47ce", 
X"47c4", X"47b9", X"47af", X"47a5", X"479a", X"4790", X"4785", X"477b", 
X"4770", X"4766", X"475c", X"4751", X"4747", X"473c", X"4732", X"4727", 
X"471d", X"4712", X"4708", X"46fe", X"46f3", X"46e9", X"46de", X"46d4", 
X"46c9", X"46bf", X"46b4", X"46aa", X"469f", X"4695", X"468a", X"4680", 
X"4675", X"466b", X"4660", X"4656", X"464b", X"4641", X"4636", X"462c", 
X"4621", X"4617", X"460c", X"4602", X"45f7", X"45ed", X"45e2", X"45d8", 
X"45cd", X"45c3", X"45b8", X"45ae", X"45a3", X"4599", X"458e", X"4583", 
X"4579", X"456e", X"4564", X"4559", X"454f", X"4544", X"4539", X"452f", 
X"4524", X"451a", X"450f", X"4505", X"44fa", X"44ef", X"44e5", X"44da", 
X"44d0", X"44c5", X"44ba", X"44b0", X"44a5", X"449b", X"4490", X"4485", 
X"447b", X"4470", X"4466", X"445b", X"4450", X"4446", X"443b", X"4430", 
X"4426", X"441b", X"4411", X"4406", X"43fb", X"43f1", X"43e6", X"43db", 
X"43d1", X"43c6", X"43bb", X"43b1", X"43a6", X"439b", X"4391", X"4386", 
X"437b", X"4371", X"4366", X"435b", X"4351", X"4346", X"433b", X"4330", 
X"4326", X"431b", X"4310", X"4306", X"42fb", X"42f0", X"42e6", X"42db", 
X"42d0", X"42c5", X"42bb", X"42b0", X"42a5", X"429a", X"4290", X"4285", 
X"427a", X"4270", X"4265", X"425a", X"424f", X"4245", X"423a", X"422f", 
X"4224", X"421a", X"420f", X"4204", X"41f9", X"41ee", X"41e4", X"41d9", 
X"41ce", X"41c3", X"41b9", X"41ae", X"41a3", X"4198", X"418d", X"4183", 
X"4178", X"416d", X"4162", X"4157", X"414d", X"4142", X"4137", X"412c", 
X"4121", X"4117", X"410c", X"4101", X"40f6", X"40eb", X"40e0", X"40d6", 
X"40cb", X"40c0", X"40b5", X"40aa", X"409f", X"4095", X"408a", X"407f", 
X"4074", X"4069", X"405e", X"4053", X"4048", X"403e", X"4033", X"4028", 
X"401d", X"4012", X"4007", X"3ffc", X"3ff1", X"3fe7", X"3fdc", X"3fd1", 
X"3fc6", X"3fbb", X"3fb0", X"3fa5", X"3f9a", X"3f8f", X"3f85", X"3f7a", 
X"3f6f", X"3f64", X"3f59", X"3f4e", X"3f43", X"3f38", X"3f2d", X"3f22", 
X"3f17", X"3f0c", X"3f01", X"3ef6", X"3eec", X"3ee1", X"3ed6", X"3ecb", 
X"3ec0", X"3eb5", X"3eaa", X"3e9f", X"3e94", X"3e89", X"3e7e", X"3e73", 
X"3e68", X"3e5d", X"3e52", X"3e47", X"3e3c", X"3e31", X"3e26", X"3e1b", 
X"3e10", X"3e05", X"3dfa", X"3def", X"3de4", X"3dd9", X"3dce", X"3dc3", 
X"3db8", X"3dad", X"3da2", X"3d97", X"3d8c", X"3d81", X"3d76", X"3d6b", 
X"3d60", X"3d55", X"3d4a", X"3d3f", X"3d34", X"3d29", X"3d1e", X"3d13", 
X"3d08", X"3cfd", X"3cf2", X"3ce7", X"3cdc", X"3cd0", X"3cc5", X"3cba", 
X"3caf", X"3ca4", X"3c99", X"3c8e", X"3c83", X"3c78", X"3c6d", X"3c62", 
X"3c57", X"3c4c", X"3c41", X"3c35", X"3c2a", X"3c1f", X"3c14", X"3c09", 
X"3bfe", X"3bf3", X"3be8", X"3bdd", X"3bd2", X"3bc6", X"3bbb", X"3bb0", 
X"3ba5", X"3b9a", X"3b8f", X"3b84", X"3b79", X"3b6d", X"3b62", X"3b57", 
X"3b4c", X"3b41", X"3b36", X"3b2b", X"3b20", X"3b14", X"3b09", X"3afe", 
X"3af3", X"3ae8", X"3add", X"3ad1", X"3ac6", X"3abb", X"3ab0", X"3aa5", 
X"3a9a", X"3a8e", X"3a83", X"3a78", X"3a6d", X"3a62", X"3a57", X"3a4b", 
X"3a40", X"3a35", X"3a2a", X"3a1f", X"3a13", X"3a08", X"39fd", X"39f2", 
X"39e7", X"39db", X"39d0", X"39c5", X"39ba", X"39af", X"39a3", X"3998", 
X"398d", X"3982", X"3976", X"396b", X"3960", X"3955", X"3949", X"393e", 
X"3933", X"3928", X"391d", X"3911", X"3906", X"38fb", X"38f0", X"38e4", 
X"38d9", X"38ce", X"38c2", X"38b7", X"38ac", X"38a1", X"3895", X"388a", 
X"387f", X"3874", X"3868", X"385d", X"3852", X"3846", X"383b", X"3830", 
X"3825", X"3819", X"380e", X"3803", X"37f7", X"37ec", X"37e1", X"37d5", 
X"37ca", X"37bf", X"37b4", X"37a8", X"379d", X"3792", X"3786", X"377b", 
X"3770", X"3764", X"3759", X"374e", X"3742", X"3737", X"372c", X"3720", 
X"3715", X"370a", X"36fe", X"36f3", X"36e8", X"36dc", X"36d1", X"36c5", 
X"36ba", X"36af", X"36a3", X"3698", X"368d", X"3681", X"3676", X"366b", 
X"365f", X"3654", X"3648", X"363d", X"3632", X"3626", X"361b", X"360f", 
X"3604", X"35f9", X"35ed", X"35e2", X"35d7", X"35cb", X"35c0", X"35b4", 
X"35a9", X"359d", X"3592", X"3587", X"357b", X"3570", X"3564", X"3559", 
X"354e", X"3542", X"3537", X"352b", X"3520", X"3514", X"3509", X"34fe", 
X"34f2", X"34e7", X"34db", X"34d0", X"34c4", X"34b9", X"34ad", X"34a2", 
X"3497", X"348b", X"3480", X"3474", X"3469", X"345d", X"3452", X"3446", 
X"343b", X"342f", X"3424", X"3418", X"340d", X"3401", X"33f6", X"33ea", 
X"33df", X"33d3", X"33c8", X"33bc", X"33b1", X"33a5", X"339a", X"338e", 
X"3383", X"3377", X"336c", X"3360", X"3355", X"3349", X"333e", X"3332", 
X"3327", X"331b", X"3310", X"3304", X"32f9", X"32ed", X"32e2", X"32d6", 
X"32cb", X"32bf", X"32b4", X"32a8", X"329d", X"3291", X"3285", X"327a", 
X"326e", X"3263", X"3257", X"324c", X"3240", X"3235", X"3229", X"321d", 
X"3212", X"3206", X"31fb", X"31ef", X"31e4", X"31d8", X"31cc", X"31c1", 
X"31b5", X"31aa", X"319e", X"3193", X"3187", X"317b", X"3170", X"3164", 
X"3159", X"314d", X"3141", X"3136", X"312a", X"311f", X"3113", X"3107", 
X"30fc", X"30f0", X"30e5", X"30d9", X"30cd", X"30c2", X"30b6", X"30aa", 
X"309f", X"3093", X"3088", X"307c", X"3070", X"3065", X"3059", X"304d", 
X"3042", X"3036", X"302a", X"301f", X"3013", X"3008", X"2ffc", X"2ff0", 
X"2fe5", X"2fd9", X"2fcd", X"2fc2", X"2fb6", X"2faa", X"2f9f", X"2f93", 
X"2f87", X"2f7c", X"2f70", X"2f64", X"2f59", X"2f4d", X"2f41", X"2f36", 
X"2f2a", X"2f1e", X"2f13", X"2f07", X"2efb", X"2eef", X"2ee4", X"2ed8", 
X"2ecc", X"2ec1", X"2eb5", X"2ea9", X"2e9e", X"2e92", X"2e86", X"2e7a", 
X"2e6f", X"2e63", X"2e57", X"2e4c", X"2e40", X"2e34", X"2e28", X"2e1d", 
X"2e11", X"2e05", X"2dfa", X"2dee", X"2de2", X"2dd6", X"2dcb", X"2dbf", 
X"2db3", X"2da7", X"2d9c", X"2d90", X"2d84", X"2d78", X"2d6d", X"2d61", 
X"2d55", X"2d49", X"2d3e", X"2d32", X"2d26", X"2d1a", X"2d0f", X"2d03", 
X"2cf7", X"2ceb", X"2ce0", X"2cd4", X"2cc8", X"2cbc", X"2cb1", X"2ca5", 
X"2c99", X"2c8d", X"2c81", X"2c76", X"2c6a", X"2c5e", X"2c52", X"2c46", 
X"2c3b", X"2c2f", X"2c23", X"2c17", X"2c0c", X"2c00", X"2bf4", X"2be8", 
X"2bdc", X"2bd0", X"2bc5", X"2bb9", X"2bad", X"2ba1", X"2b95", X"2b8a", 
X"2b7e", X"2b72", X"2b66", X"2b5a", X"2b4f", X"2b43", X"2b37", X"2b2b", 
X"2b1f", X"2b13", X"2b08", X"2afc", X"2af0", X"2ae4", X"2ad8", X"2acc", 
X"2ac1", X"2ab5", X"2aa9", X"2a9d", X"2a91", X"2a85", X"2a79", X"2a6e", 
X"2a62", X"2a56", X"2a4a", X"2a3e", X"2a32", X"2a26", X"2a1b", X"2a0f", 
X"2a03", X"29f7", X"29eb", X"29df", X"29d3", X"29c7", X"29bc", X"29b0", 
X"29a4", X"2998", X"298c", X"2980", X"2974", X"2968", X"295c", X"2951", 
X"2945", X"2939", X"292d", X"2921", X"2915", X"2909", X"28fd", X"28f1", 
X"28e5", X"28da", X"28ce", X"28c2", X"28b6", X"28aa", X"289e", X"2892", 
X"2886", X"287a", X"286e", X"2862", X"2856", X"284b", X"283f", X"2833", 
X"2827", X"281b", X"280f", X"2803", X"27f7", X"27eb", X"27df", X"27d3", 
X"27c7", X"27bb", X"27af", X"27a3", X"2797", X"278b", X"2780", X"2774", 
X"2768", X"275c", X"2750", X"2744", X"2738", X"272c", X"2720", X"2714", 
X"2708", X"26fc", X"26f0", X"26e4", X"26d8", X"26cc", X"26c0", X"26b4", 
X"26a8", X"269c", X"2690", X"2684", X"2678", X"266c", X"2660", X"2654", 
X"2648", X"263c", X"2630", X"2624", X"2618", X"260c", X"2600", X"25f4", 
X"25e8", X"25dc", X"25d0", X"25c4", X"25b8", X"25ac", X"25a0", X"2594", 
X"2588", X"257c", X"2570", X"2564", X"2558", X"254c", X"2540", X"2534", 
X"2528", X"251c", X"2510", X"2504", X"24f8", X"24ec", X"24e0", X"24d4", 
X"24c8", X"24bc", X"24b0", X"24a4", X"2498", X"248c", X"2480", X"2474", 
X"2467", X"245b", X"244f", X"2443", X"2437", X"242b", X"241f", X"2413", 
X"2407", X"23fb", X"23ef", X"23e3", X"23d7", X"23cb", X"23bf", X"23b3", 
X"23a7", X"239a", X"238e", X"2382", X"2376", X"236a", X"235e", X"2352", 
X"2346", X"233a", X"232e", X"2322", X"2316", X"230a", X"22fd", X"22f1", 
X"22e5", X"22d9", X"22cd", X"22c1", X"22b5", X"22a9", X"229d", X"2291", 
X"2284", X"2278", X"226c", X"2260", X"2254", X"2248", X"223c", X"2230", 
X"2224", X"2218", X"220b", X"21ff", X"21f3", X"21e7", X"21db", X"21cf", 
X"21c3", X"21b7", X"21aa", X"219e", X"2192", X"2186", X"217a", X"216e", 
X"2162", X"2156", X"2149", X"213d", X"2131", X"2125", X"2119", X"210d", 
X"2101", X"20f4", X"20e8", X"20dc", X"20d0", X"20c4", X"20b8", X"20ac", 
X"209f", X"2093", X"2087", X"207b", X"206f", X"2063", X"2057", X"204a", 
X"203e", X"2032", X"2026", X"201a", X"200e", X"2001", X"1ff5", X"1fe9", 
X"1fdd", X"1fd1", X"1fc5", X"1fb8", X"1fac", X"1fa0", X"1f94", X"1f88", 
X"1f7b", X"1f6f", X"1f63", X"1f57", X"1f4b", X"1f3f", X"1f32", X"1f26", 
X"1f1a", X"1f0e", X"1f02", X"1ef5", X"1ee9", X"1edd", X"1ed1", X"1ec5", 
X"1eb8", X"1eac", X"1ea0", X"1e94", X"1e88", X"1e7b", X"1e6f", X"1e63", 
X"1e57", X"1e4b", X"1e3e", X"1e32", X"1e26", X"1e1a", X"1e0e", X"1e01", 
X"1df5", X"1de9", X"1ddd", X"1dd0", X"1dc4", X"1db8", X"1dac", X"1da0", 
X"1d93", X"1d87", X"1d7b", X"1d6f", X"1d62", X"1d56", X"1d4a", X"1d3e", 
X"1d31", X"1d25", X"1d19", X"1d0d", X"1d01", X"1cf4", X"1ce8", X"1cdc", 
X"1cd0", X"1cc3", X"1cb7", X"1cab", X"1c9f", X"1c92", X"1c86", X"1c7a", 
X"1c6e", X"1c61", X"1c55", X"1c49", X"1c3d", X"1c30", X"1c24", X"1c18", 
X"1c0c", X"1bff", X"1bf3", X"1be7", X"1bda", X"1bce", X"1bc2", X"1bb6", 
X"1ba9", X"1b9d", X"1b91", X"1b85", X"1b78", X"1b6c", X"1b60", X"1b53", 
X"1b47", X"1b3b", X"1b2f", X"1b22", X"1b16", X"1b0a", X"1afe", X"1af1", 
X"1ae5", X"1ad9", X"1acc", X"1ac0", X"1ab4", X"1aa8", X"1a9b", X"1a8f", 
X"1a83", X"1a76", X"1a6a", X"1a5e", X"1a51", X"1a45", X"1a39", X"1a2d", 
X"1a20", X"1a14", X"1a08", X"19fb", X"19ef", X"19e3", X"19d6", X"19ca", 
X"19be", X"19b1", X"19a5", X"1999", X"198d", X"1980", X"1974", X"1968", 
X"195b", X"194f", X"1943", X"1936", X"192a", X"191e", X"1911", X"1905", 
X"18f9", X"18ec", X"18e0", X"18d4", X"18c7", X"18bb", X"18af", X"18a2", 
X"1896", X"188a", X"187d", X"1871", X"1865", X"1858", X"184c", X"1840", 
X"1833", X"1827", X"181b", X"180e", X"1802", X"17f6", X"17e9", X"17dd", 
X"17d1", X"17c4", X"17b8", X"17ac", X"179f", X"1793", X"1787", X"177a", 
X"176e", X"1761", X"1755", X"1749", X"173c", X"1730", X"1724", X"1717", 
X"170b", X"16ff", X"16f2", X"16e6", X"16da", X"16cd", X"16c1", X"16b4", 
X"16a8", X"169c", X"168f", X"1683", X"1677", X"166a", X"165e", X"1651", 
X"1645", X"1639", X"162c", X"1620", X"1614", X"1607", X"15fb", X"15ee", 
X"15e2", X"15d6", X"15c9", X"15bd", X"15b1", X"15a4", X"1598", X"158b", 
X"157f", X"1573", X"1566", X"155a", X"154d", X"1541", X"1535", X"1528", 
X"151c", X"150f", X"1503", X"14f7", X"14ea", X"14de", X"14d1", X"14c5", 
X"14b9", X"14ac", X"14a0", X"1493", X"1487", X"147b", X"146e", X"1462", 
X"1455", X"1449", X"143d", X"1430", X"1424", X"1417", X"140b", X"13ff", 
X"13f2", X"13e6", X"13d9", X"13cd", X"13c1", X"13b4", X"13a8", X"139b", 
X"138f", X"1382", X"1376", X"136a", X"135d", X"1351", X"1344", X"1338", 
X"132b", X"131f", X"1313", X"1306", X"12fa", X"12ed", X"12e1", X"12d4", 
X"12c8", X"12bc", X"12af", X"12a3", X"1296", X"128a", X"127d", X"1271", 
X"1265", X"1258", X"124c", X"123f", X"1233", X"1226", X"121a", X"120e", 
X"1201", X"11f5", X"11e8", X"11dc", X"11cf", X"11c3", X"11b6", X"11aa", 
X"119e", X"1191", X"1185", X"1178", X"116c", X"115f", X"1153", X"1146", 
X"113a", X"112d", X"1121", X"1115", X"1108", X"10fc", X"10ef", X"10e3", 
X"10d6", X"10ca", X"10bd", X"10b1", X"10a4", X"1098", X"108c", X"107f", 
X"1073", X"1066", X"105a", X"104d", X"1041", X"1034", X"1028", X"101b", 
X"100f", X"1002", X"0ff6", X"0fea", X"0fdd", X"0fd1", X"0fc4", X"0fb8", 
X"0fab", X"0f9f", X"0f92", X"0f86", X"0f79", X"0f6d", X"0f60", X"0f54", 
X"0f47", X"0f3b", X"0f2e", X"0f22", X"0f15", X"0f09", X"0efc", X"0ef0", 
X"0ee4", X"0ed7", X"0ecb", X"0ebe", X"0eb2", X"0ea5", X"0e99", X"0e8c", 
X"0e80", X"0e73", X"0e67", X"0e5a", X"0e4e", X"0e41", X"0e35", X"0e28", 
X"0e1c", X"0e0f", X"0e03", X"0df6", X"0dea", X"0ddd", X"0dd1", X"0dc4", 
X"0db8", X"0dab", X"0d9f", X"0d92", X"0d86", X"0d79", X"0d6d", X"0d60", 
X"0d54", X"0d47", X"0d3b", X"0d2e", X"0d22", X"0d15", X"0d09", X"0cfc", 
X"0cf0", X"0ce3", X"0cd7", X"0cca", X"0cbe", X"0cb1", X"0ca5", X"0c98", 
X"0c8c", X"0c7f", X"0c73", X"0c66", X"0c5a", X"0c4d", X"0c41", X"0c34", 
X"0c28", X"0c1b", X"0c0f", X"0c02", X"0bf6", X"0be9", X"0bdd", X"0bd0", 
X"0bc4", X"0bb7", X"0bab", X"0b9e", X"0b92", X"0b85", X"0b79", X"0b6c", 
X"0b60", X"0b53", X"0b47", X"0b3a", X"0b2d", X"0b21", X"0b14", X"0b08", 
X"0afb", X"0aef", X"0ae2", X"0ad6", X"0ac9", X"0abd", X"0ab0", X"0aa4", 
X"0a97", X"0a8b", X"0a7e", X"0a72", X"0a65", X"0a59", X"0a4c", X"0a40", 
X"0a33", X"0a27", X"0a1a", X"0a0d", X"0a01", X"09f4", X"09e8", X"09db", 
X"09cf", X"09c2", X"09b6", X"09a9", X"099d", X"0990", X"0984", X"0977", 
X"096b", X"095e", X"0951", X"0945", X"0938", X"092c", X"091f", X"0913", 
X"0906", X"08fa", X"08ed", X"08e1", X"08d4", X"08c8", X"08bb", X"08af", 
X"08a2", X"0895", X"0889", X"087c", X"0870", X"0863", X"0857", X"084a", 
X"083e", X"0831", X"0825", X"0818", X"080c", X"07ff", X"07f2", X"07e6", 
X"07d9", X"07cd", X"07c0", X"07b4", X"07a7", X"079b", X"078e", X"0782", 
X"0775", X"0768", X"075c", X"074f", X"0743", X"0736", X"072a", X"071d", 
X"0711", X"0704", X"06f8", X"06eb", X"06de", X"06d2", X"06c5", X"06b9", 
X"06ac", X"06a0", X"0693", X"0687", X"067a", X"066e", X"0661", X"0654", 
X"0648", X"063b", X"062f", X"0622", X"0616", X"0609", X"05fd", X"05f0", 
X"05e3", X"05d7", X"05ca", X"05be", X"05b1", X"05a5", X"0598", X"058c", 
X"057f", X"0572", X"0566", X"0559", X"054d", X"0540", X"0534", X"0527", 
X"051b", X"050e", X"0501", X"04f5", X"04e8", X"04dc", X"04cf", X"04c3", 
X"04b6", X"04aa", X"049d", X"0490", X"0484", X"0477", X"046b", X"045e", 
X"0452", X"0445", X"0439", X"042c", X"041f", X"0413", X"0406", X"03fa", 
X"03ed", X"03e1", X"03d4", X"03c7", X"03bb", X"03ae", X"03a2", X"0395", 
X"0389", X"037c", X"0370", X"0363", X"0356", X"034a", X"033d", X"0331", 
X"0324", X"0318", X"030b", X"02fe", X"02f2", X"02e5", X"02d9", X"02cc", 
X"02c0", X"02b3", X"02a7", X"029a", X"028d", X"0281", X"0274", X"0268", 
X"025b", X"024f", X"0242", X"0235", X"0229", X"021c", X"0210", X"0203", 
X"01f7", X"01ea", X"01de", X"01d1", X"01c4", X"01b8", X"01ab", X"019f", 
X"0192", X"0186", X"0179", X"016c", X"0160", X"0153", X"0147", X"013a", 
X"012e", X"0121", X"0114", X"0108", X"00fb", X"00ef", X"00e2", X"00d6", 
X"00c9", X"00bc", X"00b0", X"00a3", X"0097", X"008a", X"007e", X"0071", 
X"0065", X"0058", X"004b", X"003f", X"0032", X"0026", X"0019", X"000d", 
X"0000", X"fff3", X"ffe7", X"ffda", X"ffce", X"ffc1", X"ffb5", X"ffa8", 
X"ff9b", X"ff8f", X"ff82", X"ff76", X"ff69", X"ff5d", X"ff50", X"ff44", 
X"ff37", X"ff2a", X"ff1e", X"ff11", X"ff05", X"fef8", X"feec", X"fedf", 
X"fed2", X"fec6", X"feb9", X"fead", X"fea0", X"fe94", X"fe87", X"fe7a", 
X"fe6e", X"fe61", X"fe55", X"fe48", X"fe3c", X"fe2f", X"fe22", X"fe16", 
X"fe09", X"fdfd", X"fdf0", X"fde4", X"fdd7", X"fdcb", X"fdbe", X"fdb1", 
X"fda5", X"fd98", X"fd8c", X"fd7f", X"fd73", X"fd66", X"fd59", X"fd4d", 
X"fd40", X"fd34", X"fd27", X"fd1b", X"fd0e", X"fd02", X"fcf5", X"fce8", 
X"fcdc", X"fccf", X"fcc3", X"fcb6", X"fcaa", X"fc9d", X"fc90", X"fc84", 
X"fc77", X"fc6b", X"fc5e", X"fc52", X"fc45", X"fc39", X"fc2c", X"fc1f", 
X"fc13", X"fc06", X"fbfa", X"fbed", X"fbe1", X"fbd4", X"fbc7", X"fbbb", 
X"fbae", X"fba2", X"fb95", X"fb89", X"fb7c", X"fb70", X"fb63", X"fb56", 
X"fb4a", X"fb3d", X"fb31", X"fb24", X"fb18", X"fb0b", X"faff", X"faf2", 
X"fae5", X"fad9", X"facc", X"fac0", X"fab3", X"faa7", X"fa9a", X"fa8e", 
X"fa81", X"fa74", X"fa68", X"fa5b", X"fa4f", X"fa42", X"fa36", X"fa29", 
X"fa1d", X"fa10", X"fa03", X"f9f7", X"f9ea", X"f9de", X"f9d1", X"f9c5", 
X"f9b8", X"f9ac", X"f99f", X"f992", X"f986", X"f979", X"f96d", X"f960", 
X"f954", X"f947", X"f93b", X"f92e", X"f922", X"f915", X"f908", X"f8fc", 
X"f8ef", X"f8e3", X"f8d6", X"f8ca", X"f8bd", X"f8b1", X"f8a4", X"f898", 
X"f88b", X"f87e", X"f872", X"f865", X"f859", X"f84c", X"f840", X"f833", 
X"f827", X"f81a", X"f80e", X"f801", X"f7f4", X"f7e8", X"f7db", X"f7cf", 
X"f7c2", X"f7b6", X"f7a9", X"f79d", X"f790", X"f784", X"f777", X"f76b", 
X"f75e", X"f751", X"f745", X"f738", X"f72c", X"f71f", X"f713", X"f706", 
X"f6fa", X"f6ed", X"f6e1", X"f6d4", X"f6c8", X"f6bb", X"f6af", X"f6a2", 
X"f695", X"f689", X"f67c", X"f670", X"f663", X"f657", X"f64a", X"f63e", 
X"f631", X"f625", X"f618", X"f60c", X"f5ff", X"f5f3", X"f5e6", X"f5d9", 
X"f5cd", X"f5c0", X"f5b4", X"f5a7", X"f59b", X"f58e", X"f582", X"f575", 
X"f569", X"f55c", X"f550", X"f543", X"f537", X"f52a", X"f51e", X"f511", 
X"f505", X"f4f8", X"f4ec", X"f4df", X"f4d3", X"f4c6", X"f4b9", X"f4ad", 
X"f4a0", X"f494", X"f487", X"f47b", X"f46e", X"f462", X"f455", X"f449", 
X"f43c", X"f430", X"f423", X"f417", X"f40a", X"f3fe", X"f3f1", X"f3e5", 
X"f3d8", X"f3cc", X"f3bf", X"f3b3", X"f3a6", X"f39a", X"f38d", X"f381", 
X"f374", X"f368", X"f35b", X"f34f", X"f342", X"f336", X"f329", X"f31d", 
X"f310", X"f304", X"f2f7", X"f2eb", X"f2de", X"f2d2", X"f2c5", X"f2b9", 
X"f2ac", X"f2a0", X"f293", X"f287", X"f27a", X"f26e", X"f261", X"f255", 
X"f248", X"f23c", X"f22f", X"f223", X"f216", X"f20a", X"f1fd", X"f1f1", 
X"f1e4", X"f1d8", X"f1cb", X"f1bf", X"f1b2", X"f1a6", X"f199", X"f18d", 
X"f180", X"f174", X"f167", X"f15b", X"f14e", X"f142", X"f135", X"f129", 
X"f11c", X"f110", X"f104", X"f0f7", X"f0eb", X"f0de", X"f0d2", X"f0c5", 
X"f0b9", X"f0ac", X"f0a0", X"f093", X"f087", X"f07a", X"f06e", X"f061", 
X"f055", X"f048", X"f03c", X"f02f", X"f023", X"f016", X"f00a", X"effe", 
X"eff1", X"efe5", X"efd8", X"efcc", X"efbf", X"efb3", X"efa6", X"ef9a", 
X"ef8d", X"ef81", X"ef74", X"ef68", X"ef5c", X"ef4f", X"ef43", X"ef36", 
X"ef2a", X"ef1d", X"ef11", X"ef04", X"eef8", X"eeeb", X"eedf", X"eed3", 
X"eec6", X"eeba", X"eead", X"eea1", X"ee94", X"ee88", X"ee7b", X"ee6f", 
X"ee62", X"ee56", X"ee4a", X"ee3d", X"ee31", X"ee24", X"ee18", X"ee0b", 
X"edff", X"edf2", X"ede6", X"edda", X"edcd", X"edc1", X"edb4", X"eda8", 
X"ed9b", X"ed8f", X"ed83", X"ed76", X"ed6a", X"ed5d", X"ed51", X"ed44", 
X"ed38", X"ed2c", X"ed1f", X"ed13", X"ed06", X"ecfa", X"eced", X"ece1", 
X"ecd5", X"ecc8", X"ecbc", X"ecaf", X"eca3", X"ec96", X"ec8a", X"ec7e", 
X"ec71", X"ec65", X"ec58", X"ec4c", X"ec3f", X"ec33", X"ec27", X"ec1a", 
X"ec0e", X"ec01", X"ebf5", X"ebe9", X"ebdc", X"ebd0", X"ebc3", X"ebb7", 
X"ebab", X"eb9e", X"eb92", X"eb85", X"eb79", X"eb6d", X"eb60", X"eb54", 
X"eb47", X"eb3b", X"eb2f", X"eb22", X"eb16", X"eb09", X"eafd", X"eaf1", 
X"eae4", X"ead8", X"eacb", X"eabf", X"eab3", X"eaa6", X"ea9a", X"ea8d", 
X"ea81", X"ea75", X"ea68", X"ea5c", X"ea4f", X"ea43", X"ea37", X"ea2a", 
X"ea1e", X"ea12", X"ea05", X"e9f9", X"e9ec", X"e9e0", X"e9d4", X"e9c7", 
X"e9bb", X"e9af", X"e9a2", X"e996", X"e989", X"e97d", X"e971", X"e964", 
X"e958", X"e94c", X"e93f", X"e933", X"e926", X"e91a", X"e90e", X"e901", 
X"e8f5", X"e8e9", X"e8dc", X"e8d0", X"e8c4", X"e8b7", X"e8ab", X"e89f", 
X"e892", X"e886", X"e879", X"e86d", X"e861", X"e854", X"e848", X"e83c", 
X"e82f", X"e823", X"e817", X"e80a", X"e7fe", X"e7f2", X"e7e5", X"e7d9", 
X"e7cd", X"e7c0", X"e7b4", X"e7a8", X"e79b", X"e78f", X"e783", X"e776", 
X"e76a", X"e75e", X"e751", X"e745", X"e739", X"e72c", X"e720", X"e714", 
X"e707", X"e6fb", X"e6ef", X"e6e2", X"e6d6", X"e6ca", X"e6bd", X"e6b1", 
X"e6a5", X"e698", X"e68c", X"e680", X"e673", X"e667", X"e65b", X"e64f", 
X"e642", X"e636", X"e62a", X"e61d", X"e611", X"e605", X"e5f8", X"e5ec", 
X"e5e0", X"e5d3", X"e5c7", X"e5bb", X"e5af", X"e5a2", X"e596", X"e58a", 
X"e57d", X"e571", X"e565", X"e558", X"e54c", X"e540", X"e534", X"e527", 
X"e51b", X"e50f", X"e502", X"e4f6", X"e4ea", X"e4de", X"e4d1", X"e4c5", 
X"e4b9", X"e4ad", X"e4a0", X"e494", X"e488", X"e47b", X"e46f", X"e463", 
X"e457", X"e44a", X"e43e", X"e432", X"e426", X"e419", X"e40d", X"e401", 
X"e3f4", X"e3e8", X"e3dc", X"e3d0", X"e3c3", X"e3b7", X"e3ab", X"e39f", 
X"e392", X"e386", X"e37a", X"e36e", X"e361", X"e355", X"e349", X"e33d", 
X"e330", X"e324", X"e318", X"e30c", X"e2ff", X"e2f3", X"e2e7", X"e2db", 
X"e2cf", X"e2c2", X"e2b6", X"e2aa", X"e29e", X"e291", X"e285", X"e279", 
X"e26d", X"e260", X"e254", X"e248", X"e23c", X"e230", X"e223", X"e217", 
X"e20b", X"e1ff", X"e1f2", X"e1e6", X"e1da", X"e1ce", X"e1c2", X"e1b5", 
X"e1a9", X"e19d", X"e191", X"e185", X"e178", X"e16c", X"e160", X"e154", 
X"e148", X"e13b", X"e12f", X"e123", X"e117", X"e10b", X"e0fe", X"e0f2", 
X"e0e6", X"e0da", X"e0ce", X"e0c1", X"e0b5", X"e0a9", X"e09d", X"e091", 
X"e085", X"e078", X"e06c", X"e060", X"e054", X"e048", X"e03b", X"e02f", 
X"e023", X"e017", X"e00b", X"dfff", X"dff2", X"dfe6", X"dfda", X"dfce", 
X"dfc2", X"dfb6", X"dfa9", X"df9d", X"df91", X"df85", X"df79", X"df6d", 
X"df61", X"df54", X"df48", X"df3c", X"df30", X"df24", X"df18", X"df0c", 
X"deff", X"def3", X"dee7", X"dedb", X"decf", X"dec3", X"deb7", X"deaa", 
X"de9e", X"de92", X"de86", X"de7a", X"de6e", X"de62", X"de56", X"de49", 
X"de3d", X"de31", X"de25", X"de19", X"de0d", X"de01", X"ddf5", X"dde8", 
X"dddc", X"ddd0", X"ddc4", X"ddb8", X"ddac", X"dda0", X"dd94", X"dd88", 
X"dd7c", X"dd6f", X"dd63", X"dd57", X"dd4b", X"dd3f", X"dd33", X"dd27", 
X"dd1b", X"dd0f", X"dd03", X"dcf6", X"dcea", X"dcde", X"dcd2", X"dcc6", 
X"dcba", X"dcae", X"dca2", X"dc96", X"dc8a", X"dc7e", X"dc72", X"dc66", 
X"dc59", X"dc4d", X"dc41", X"dc35", X"dc29", X"dc1d", X"dc11", X"dc05", 
X"dbf9", X"dbed", X"dbe1", X"dbd5", X"dbc9", X"dbbd", X"dbb1", X"dba5", 
X"db99", X"db8c", X"db80", X"db74", X"db68", X"db5c", X"db50", X"db44", 
X"db38", X"db2c", X"db20", X"db14", X"db08", X"dafc", X"daf0", X"dae4", 
X"dad8", X"dacc", X"dac0", X"dab4", X"daa8", X"da9c", X"da90", X"da84", 
X"da78", X"da6c", X"da60", X"da54", X"da48", X"da3c", X"da30", X"da24", 
X"da18", X"da0c", X"da00", X"d9f4", X"d9e8", X"d9dc", X"d9d0", X"d9c4", 
X"d9b8", X"d9ac", X"d9a0", X"d994", X"d988", X"d97c", X"d970", X"d964", 
X"d958", X"d94c", X"d940", X"d934", X"d928", X"d91c", X"d910", X"d904", 
X"d8f8", X"d8ec", X"d8e0", X"d8d4", X"d8c8", X"d8bc", X"d8b0", X"d8a4", 
X"d898", X"d88c", X"d880", X"d875", X"d869", X"d85d", X"d851", X"d845", 
X"d839", X"d82d", X"d821", X"d815", X"d809", X"d7fd", X"d7f1", X"d7e5", 
X"d7d9", X"d7cd", X"d7c1", X"d7b5", X"d7aa", X"d79e", X"d792", X"d786", 
X"d77a", X"d76e", X"d762", X"d756", X"d74a", X"d73e", X"d732", X"d726", 
X"d71b", X"d70f", X"d703", X"d6f7", X"d6eb", X"d6df", X"d6d3", X"d6c7", 
X"d6bb", X"d6af", X"d6a4", X"d698", X"d68c", X"d680", X"d674", X"d668", 
X"d65c", X"d650", X"d644", X"d639", X"d62d", X"d621", X"d615", X"d609", 
X"d5fd", X"d5f1", X"d5e5", X"d5da", X"d5ce", X"d5c2", X"d5b6", X"d5aa", 
X"d59e", X"d592", X"d587", X"d57b", X"d56f", X"d563", X"d557", X"d54b", 
X"d53f", X"d534", X"d528", X"d51c", X"d510", X"d504", X"d4f8", X"d4ed", 
X"d4e1", X"d4d5", X"d4c9", X"d4bd", X"d4b1", X"d4a6", X"d49a", X"d48e", 
X"d482", X"d476", X"d46b", X"d45f", X"d453", X"d447", X"d43b", X"d430", 
X"d424", X"d418", X"d40c", X"d400", X"d3f4", X"d3e9", X"d3dd", X"d3d1", 
X"d3c5", X"d3ba", X"d3ae", X"d3a2", X"d396", X"d38a", X"d37f", X"d373", 
X"d367", X"d35b", X"d34f", X"d344", X"d338", X"d32c", X"d320", X"d315", 
X"d309", X"d2fd", X"d2f1", X"d2e6", X"d2da", X"d2ce", X"d2c2", X"d2b7", 
X"d2ab", X"d29f", X"d293", X"d288", X"d27c", X"d270", X"d264", X"d259", 
X"d24d", X"d241", X"d235", X"d22a", X"d21e", X"d212", X"d206", X"d1fb", 
X"d1ef", X"d1e3", X"d1d8", X"d1cc", X"d1c0", X"d1b4", X"d1a9", X"d19d", 
X"d191", X"d186", X"d17a", X"d16e", X"d162", X"d157", X"d14b", X"d13f", 
X"d134", X"d128", X"d11c", X"d111", X"d105", X"d0f9", X"d0ed", X"d0e2", 
X"d0d6", X"d0ca", X"d0bf", X"d0b3", X"d0a7", X"d09c", X"d090", X"d084", 
X"d079", X"d06d", X"d061", X"d056", X"d04a", X"d03e", X"d033", X"d027", 
X"d01b", X"d010", X"d004", X"cff8", X"cfed", X"cfe1", X"cfd6", X"cfca", 
X"cfbe", X"cfb3", X"cfa7", X"cf9b", X"cf90", X"cf84", X"cf78", X"cf6d", 
X"cf61", X"cf56", X"cf4a", X"cf3e", X"cf33", X"cf27", X"cf1b", X"cf10", 
X"cf04", X"cef9", X"ceed", X"cee1", X"ced6", X"ceca", X"cebf", X"ceb3", 
X"cea7", X"ce9c", X"ce90", X"ce85", X"ce79", X"ce6d", X"ce62", X"ce56", 
X"ce4b", X"ce3f", X"ce34", X"ce28", X"ce1c", X"ce11", X"ce05", X"cdfa", 
X"cdee", X"cde3", X"cdd7", X"cdcb", X"cdc0", X"cdb4", X"cda9", X"cd9d", 
X"cd92", X"cd86", X"cd7b", X"cd6f", X"cd63", X"cd58", X"cd4c", X"cd41", 
X"cd35", X"cd2a", X"cd1e", X"cd13", X"cd07", X"ccfc", X"ccf0", X"cce5", 
X"ccd9", X"ccce", X"ccc2", X"ccb7", X"ccab", X"cca0", X"cc94", X"cc89", 
X"cc7d", X"cc72", X"cc66", X"cc5b", X"cc4f", X"cc44", X"cc38", X"cc2d", 
X"cc21", X"cc16", X"cc0a", X"cbff", X"cbf3", X"cbe8", X"cbdc", X"cbd1", 
X"cbc5", X"cbba", X"cbae", X"cba3", X"cb97", X"cb8c", X"cb80", X"cb75", 
X"cb69", X"cb5e", X"cb53", X"cb47", X"cb3c", X"cb30", X"cb25", X"cb19", 
X"cb0e", X"cb02", X"caf7", X"caec", X"cae0", X"cad5", X"cac9", X"cabe", 
X"cab2", X"caa7", X"ca9c", X"ca90", X"ca85", X"ca79", X"ca6e", X"ca63", 
X"ca57", X"ca4c", X"ca40", X"ca35", X"ca29", X"ca1e", X"ca13", X"ca07", 
X"c9fc", X"c9f1", X"c9e5", X"c9da", X"c9ce", X"c9c3", X"c9b8", X"c9ac", 
X"c9a1", X"c995", X"c98a", X"c97f", X"c973", X"c968", X"c95d", X"c951", 
X"c946", X"c93b", X"c92f", X"c924", X"c918", X"c90d", X"c902", X"c8f6", 
X"c8eb", X"c8e0", X"c8d4", X"c8c9", X"c8be", X"c8b2", X"c8a7", X"c89c", 
X"c890", X"c885", X"c87a", X"c86e", X"c863", X"c858", X"c84c", X"c841", 
X"c836", X"c82b", X"c81f", X"c814", X"c809", X"c7fd", X"c7f2", X"c7e7", 
X"c7db", X"c7d0", X"c7c5", X"c7ba", X"c7ae", X"c7a3", X"c798", X"c78c", 
X"c781", X"c776", X"c76b", X"c75f", X"c754", X"c749", X"c73e", X"c732", 
X"c727", X"c71c", X"c710", X"c705", X"c6fa", X"c6ef", X"c6e3", X"c6d8", 
X"c6cd", X"c6c2", X"c6b7", X"c6ab", X"c6a0", X"c695", X"c68a", X"c67e", 
X"c673", X"c668", X"c65d", X"c651", X"c646", X"c63b", X"c630", X"c625", 
X"c619", X"c60e", X"c603", X"c5f8", X"c5ed", X"c5e1", X"c5d6", X"c5cb", 
X"c5c0", X"c5b5", X"c5a9", X"c59e", X"c593", X"c588", X"c57d", X"c572", 
X"c566", X"c55b", X"c550", X"c545", X"c53a", X"c52f", X"c523", X"c518", 
X"c50d", X"c502", X"c4f7", X"c4ec", X"c4e0", X"c4d5", X"c4ca", X"c4bf", 
X"c4b4", X"c4a9", X"c49e", X"c493", X"c487", X"c47c", X"c471", X"c466", 
X"c45b", X"c450", X"c445", X"c43a", X"c42e", X"c423", X"c418", X"c40d", 
X"c402", X"c3f7", X"c3ec", X"c3e1", X"c3d6", X"c3cb", X"c3bf", X"c3b4", 
X"c3a9", X"c39e", X"c393", X"c388", X"c37d", X"c372", X"c367", X"c35c", 
X"c351", X"c346", X"c33b", X"c330", X"c324", X"c319", X"c30e", X"c303", 
X"c2f8", X"c2ed", X"c2e2", X"c2d7", X"c2cc", X"c2c1", X"c2b6", X"c2ab", 
X"c2a0", X"c295", X"c28a", X"c27f", X"c274", X"c269", X"c25e", X"c253", 
X"c248", X"c23d", X"c232", X"c227", X"c21c", X"c211", X"c206", X"c1fb", 
X"c1f0", X"c1e5", X"c1da", X"c1cf", X"c1c4", X"c1b9", X"c1ae", X"c1a3", 
X"c198", X"c18d", X"c182", X"c177", X"c16c", X"c161", X"c156", X"c14b", 
X"c140", X"c135", X"c12a", X"c11f", X"c114", X"c10a", X"c0ff", X"c0f4", 
X"c0e9", X"c0de", X"c0d3", X"c0c8", X"c0bd", X"c0b2", X"c0a7", X"c09c", 
X"c091", X"c086", X"c07b", X"c071", X"c066", X"c05b", X"c050", X"c045", 
X"c03a", X"c02f", X"c024", X"c019", X"c00f", X"c004", X"bff9", X"bfee", 
X"bfe3", X"bfd8", X"bfcd", X"bfc2", X"bfb8", X"bfad", X"bfa2", X"bf97", 
X"bf8c", X"bf81", X"bf76", X"bf6b", X"bf61", X"bf56", X"bf4b", X"bf40", 
X"bf35", X"bf2a", X"bf20", X"bf15", X"bf0a", X"beff", X"bef4", X"bee9", 
X"bedf", X"bed4", X"bec9", X"bebe", X"beb3", X"bea9", X"be9e", X"be93", 
X"be88", X"be7d", X"be73", X"be68", X"be5d", X"be52", X"be47", X"be3d", 
X"be32", X"be27", X"be1c", X"be12", X"be07", X"bdfc", X"bdf1", X"bde6", 
X"bddc", X"bdd1", X"bdc6", X"bdbb", X"bdb1", X"bda6", X"bd9b", X"bd90", 
X"bd86", X"bd7b", X"bd70", X"bd66", X"bd5b", X"bd50", X"bd45", X"bd3b", 
X"bd30", X"bd25", X"bd1a", X"bd10", X"bd05", X"bcfa", X"bcf0", X"bce5", 
X"bcda", X"bcd0", X"bcc5", X"bcba", X"bcaf", X"bca5", X"bc9a", X"bc8f", 
X"bc85", X"bc7a", X"bc6f", X"bc65", X"bc5a", X"bc4f", X"bc45", X"bc3a", 
X"bc2f", X"bc25", X"bc1a", X"bc0f", X"bc05", X"bbfa", X"bbef", X"bbe5", 
X"bbda", X"bbd0", X"bbc5", X"bbba", X"bbb0", X"bba5", X"bb9a", X"bb90", 
X"bb85", X"bb7b", X"bb70", X"bb65", X"bb5b", X"bb50", X"bb46", X"bb3b", 
X"bb30", X"bb26", X"bb1b", X"bb11", X"bb06", X"bafb", X"baf1", X"bae6", 
X"badc", X"bad1", X"bac7", X"babc", X"bab1", X"baa7", X"ba9c", X"ba92", 
X"ba87", X"ba7d", X"ba72", X"ba67", X"ba5d", X"ba52", X"ba48", X"ba3d", 
X"ba33", X"ba28", X"ba1e", X"ba13", X"ba09", X"b9fe", X"b9f4", X"b9e9", 
X"b9df", X"b9d4", X"b9ca", X"b9bf", X"b9b5", X"b9aa", X"b9a0", X"b995", 
X"b98b", X"b980", X"b976", X"b96b", X"b961", X"b956", X"b94c", X"b941", 
X"b937", X"b92c", X"b922", X"b917", X"b90d", X"b902", X"b8f8", X"b8ee", 
X"b8e3", X"b8d9", X"b8ce", X"b8c4", X"b8b9", X"b8af", X"b8a4", X"b89a", 
X"b890", X"b885", X"b87b", X"b870", X"b866", X"b85b", X"b851", X"b847", 
X"b83c", X"b832", X"b827", X"b81d", X"b813", X"b808", X"b7fe", X"b7f3", 
X"b7e9", X"b7df", X"b7d4", X"b7ca", X"b7c0", X"b7b5", X"b7ab", X"b7a0", 
X"b796", X"b78c", X"b781", X"b777", X"b76d", X"b762", X"b758", X"b74e", 
X"b743", X"b739", X"b72f", X"b724", X"b71a", X"b710", X"b705", X"b6fb", 
X"b6f1", X"b6e6", X"b6dc", X"b6d2", X"b6c7", X"b6bd", X"b6b3", X"b6a8", 
X"b69e", X"b694", X"b68a", X"b67f", X"b675", X"b66b", X"b660", X"b656", 
X"b64c", X"b642", X"b637", X"b62d", X"b623", X"b619", X"b60e", X"b604", 
X"b5fa", X"b5f0", X"b5e5", X"b5db", X"b5d1", X"b5c7", X"b5bc", X"b5b2", 
X"b5a8", X"b59e", X"b593", X"b589", X"b57f", X"b575", X"b56b", X"b560", 
X"b556", X"b54c", X"b542", X"b538", X"b52d", X"b523", X"b519", X"b50f", 
X"b505", X"b4fa", X"b4f0", X"b4e6", X"b4dc", X"b4d2", X"b4c8", X"b4bd", 
X"b4b3", X"b4a9", X"b49f", X"b495", X"b48b", X"b480", X"b476", X"b46c", 
X"b462", X"b458", X"b44e", X"b444", X"b439", X"b42f", X"b425", X"b41b", 
X"b411", X"b407", X"b3fd", X"b3f3", X"b3e9", X"b3de", X"b3d4", X"b3ca", 
X"b3c0", X"b3b6", X"b3ac", X"b3a2", X"b398", X"b38e", X"b384", X"b37a", 
X"b36f", X"b365", X"b35b", X"b351", X"b347", X"b33d", X"b333", X"b329", 
X"b31f", X"b315", X"b30b", X"b301", X"b2f7", X"b2ed", X"b2e3", X"b2d9", 
X"b2cf", X"b2c5", X"b2bb", X"b2b1", X"b2a7", X"b29d", X"b293", X"b289", 
X"b27f", X"b275", X"b26b", X"b261", X"b257", X"b24d", X"b243", X"b239", 
X"b22f", X"b225", X"b21b", X"b211", X"b207", X"b1fd", X"b1f3", X"b1e9", 
X"b1df", X"b1d5", X"b1cb", X"b1c1", X"b1b7", X"b1ad", X"b1a3", X"b199", 
X"b18f", X"b186", X"b17c", X"b172", X"b168", X"b15e", X"b154", X"b14a", 
X"b140", X"b136", X"b12c", X"b122", X"b118", X"b10f", X"b105", X"b0fb", 
X"b0f1", X"b0e7", X"b0dd", X"b0d3", X"b0c9", X"b0c0", X"b0b6", X"b0ac", 
X"b0a2", X"b098", X"b08e", X"b084", X"b07b", X"b071", X"b067", X"b05d", 
X"b053", X"b049", X"b040", X"b036", X"b02c", X"b022", X"b018", X"b00e", 
X"b005", X"affb", X"aff1", X"afe7", X"afdd", X"afd4", X"afca", X"afc0", 
X"afb6", X"afac", X"afa3", X"af99", X"af8f", X"af85", X"af7c", X"af72", 
X"af68", X"af5e", X"af54", X"af4b", X"af41", X"af37", X"af2d", X"af24", 
X"af1a", X"af10", X"af07", X"aefd", X"aef3", X"aee9", X"aee0", X"aed6", 
X"aecc", X"aec2", X"aeb9", X"aeaf", X"aea5", X"ae9c", X"ae92", X"ae88", 
X"ae7f", X"ae75", X"ae6b", X"ae62", X"ae58", X"ae4e", X"ae45", X"ae3b", 
X"ae31", X"ae28", X"ae1e", X"ae14", X"ae0b", X"ae01", X"adf7", X"adee", 
X"ade4", X"adda", X"add1", X"adc7", X"adbd", X"adb4", X"adaa", X"ada1", 
X"ad97", X"ad8d", X"ad84", X"ad7a", X"ad70", X"ad67", X"ad5d", X"ad54", 
X"ad4a", X"ad41", X"ad37", X"ad2d", X"ad24", X"ad1a", X"ad11", X"ad07", 
X"acfd", X"acf4", X"acea", X"ace1", X"acd7", X"acce", X"acc4", X"acbb", 
X"acb1", X"aca8", X"ac9e", X"ac94", X"ac8b", X"ac81", X"ac78", X"ac6e", 
X"ac65", X"ac5b", X"ac52", X"ac48", X"ac3f", X"ac35", X"ac2c", X"ac22", 
X"ac19", X"ac0f", X"ac06", X"abfc", X"abf3", X"abe9", X"abe0", X"abd6", 
X"abcd", X"abc4", X"abba", X"abb1", X"aba7", X"ab9e", X"ab94", X"ab8b", 
X"ab81", X"ab78", X"ab6f", X"ab65", X"ab5c", X"ab52", X"ab49", X"ab3f", 
X"ab36", X"ab2d", X"ab23", X"ab1a", X"ab10", X"ab07", X"aafe", X"aaf4", 
X"aaeb", X"aae1", X"aad8", X"aacf", X"aac5", X"aabc", X"aab2", X"aaa9", 
X"aaa0", X"aa96", X"aa8d", X"aa84", X"aa7a", X"aa71", X"aa68", X"aa5e", 
X"aa55", X"aa4c", X"aa42", X"aa39", X"aa30", X"aa26", X"aa1d", X"aa14", 
X"aa0a", X"aa01", X"a9f8", X"a9ee", X"a9e5", X"a9dc", X"a9d3", X"a9c9", 
X"a9c0", X"a9b7", X"a9ad", X"a9a4", X"a99b", X"a992", X"a988", X"a97f", 
X"a976", X"a96d", X"a963", X"a95a", X"a951", X"a948", X"a93e", X"a935", 
X"a92c", X"a923", X"a919", X"a910", X"a907", X"a8fe", X"a8f4", X"a8eb", 
X"a8e2", X"a8d9", X"a8d0", X"a8c6", X"a8bd", X"a8b4", X"a8ab", X"a8a2", 
X"a899", X"a88f", X"a886", X"a87d", X"a874", X"a86b", X"a861", X"a858", 
X"a84f", X"a846", X"a83d", X"a834", X"a82b", X"a821", X"a818", X"a80f", 
X"a806", X"a7fd", X"a7f4", X"a7eb", X"a7e2", X"a7d8", X"a7cf", X"a7c6", 
X"a7bd", X"a7b4", X"a7ab", X"a7a2", X"a799", X"a790", X"a787", X"a77e", 
X"a774", X"a76b", X"a762", X"a759", X"a750", X"a747", X"a73e", X"a735", 
X"a72c", X"a723", X"a71a", X"a711", X"a708", X"a6ff", X"a6f6", X"a6ed", 
X"a6e4", X"a6db", X"a6d2", X"a6c9", X"a6c0", X"a6b7", X"a6ae", X"a6a5", 
X"a69c", X"a693", X"a68a", X"a681", X"a678", X"a66f", X"a666", X"a65d", 
X"a654", X"a64b", X"a642", X"a639", X"a630", X"a627", X"a61e", X"a615", 
X"a60c", X"a603", X"a5fa", X"a5f1", X"a5e8", X"a5df", X"a5d7", X"a5ce", 
X"a5c5", X"a5bc", X"a5b3", X"a5aa", X"a5a1", X"a598", X"a58f", X"a586", 
X"a57e", X"a575", X"a56c", X"a563", X"a55a", X"a551", X"a548", X"a53f", 
X"a537", X"a52e", X"a525", X"a51c", X"a513", X"a50a", X"a501", X"a4f9", 
X"a4f0", X"a4e7", X"a4de", X"a4d5", X"a4cc", X"a4c4", X"a4bb", X"a4b2", 
X"a4a9", X"a4a0", X"a498", X"a48f", X"a486", X"a47d", X"a474", X"a46c", 
X"a463", X"a45a", X"a451", X"a449", X"a440", X"a437", X"a42e", X"a426", 
X"a41d", X"a414", X"a40b", X"a403", X"a3fa", X"a3f1", X"a3e8", X"a3e0", 
X"a3d7", X"a3ce", X"a3c6", X"a3bd", X"a3b4", X"a3ab", X"a3a3", X"a39a", 
X"a391", X"a389", X"a380", X"a377", X"a36f", X"a366", X"a35d", X"a355", 
X"a34c", X"a343", X"a33b", X"a332", X"a329", X"a321", X"a318", X"a30f", 
X"a307", X"a2fe", X"a2f5", X"a2ed", X"a2e4", X"a2dc", X"a2d3", X"a2ca", 
X"a2c2", X"a2b9", X"a2b0", X"a2a8", X"a29f", X"a297", X"a28e", X"a286", 
X"a27d", X"a274", X"a26c", X"a263", X"a25b", X"a252", X"a249", X"a241", 
X"a238", X"a230", X"a227", X"a21f", X"a216", X"a20e", X"a205", X"a1fd", 
X"a1f4", X"a1ec", X"a1e3", X"a1db", X"a1d2", X"a1c9", X"a1c1", X"a1b8", 
X"a1b0", X"a1a8", X"a19f", X"a197", X"a18e", X"a186", X"a17d", X"a175", 
X"a16c", X"a164", X"a15b", X"a153", X"a14a", X"a142", X"a139", X"a131", 
X"a129", X"a120", X"a118", X"a10f", X"a107", X"a0fe", X"a0f6", X"a0ee", 
X"a0e5", X"a0dd", X"a0d4", X"a0cc", X"a0c4", X"a0bb", X"a0b3", X"a0aa", 
X"a0a2", X"a09a", X"a091", X"a089", X"a080", X"a078", X"a070", X"a067", 
X"a05f", X"a057", X"a04e", X"a046", X"a03e", X"a035", X"a02d", X"a025", 
X"a01c", X"a014", X"a00c", X"a003", X"9ffb", X"9ff3", X"9fea", X"9fe2", 
X"9fda", X"9fd2", X"9fc9", X"9fc1", X"9fb9", X"9fb0", X"9fa8", X"9fa0", 
X"9f98", X"9f8f", X"9f87", X"9f7f", X"9f77", X"9f6e", X"9f66", X"9f5e", 
X"9f56", X"9f4d", X"9f45", X"9f3d", X"9f35", X"9f2c", X"9f24", X"9f1c", 
X"9f14", X"9f0c", X"9f03", X"9efb", X"9ef3", X"9eeb", X"9ee3", X"9eda", 
X"9ed2", X"9eca", X"9ec2", X"9eba", X"9eb2", X"9ea9", X"9ea1", X"9e99", 
X"9e91", X"9e89", X"9e81", X"9e78", X"9e70", X"9e68", X"9e60", X"9e58", 
X"9e50", X"9e48", X"9e40", X"9e37", X"9e2f", X"9e27", X"9e1f", X"9e17", 
X"9e0f", X"9e07", X"9dff", X"9df7", X"9def", X"9de7", X"9ddf", X"9dd6", 
X"9dce", X"9dc6", X"9dbe", X"9db6", X"9dae", X"9da6", X"9d9e", X"9d96", 
X"9d8e", X"9d86", X"9d7e", X"9d76", X"9d6e", X"9d66", X"9d5e", X"9d56", 
X"9d4e", X"9d46", X"9d3e", X"9d36", X"9d2e", X"9d26", X"9d1e", X"9d16", 
X"9d0e", X"9d06", X"9cfe", X"9cf6", X"9cee", X"9ce6", X"9cde", X"9cd6", 
X"9cce", X"9cc6", X"9cbe", X"9cb7", X"9caf", X"9ca7", X"9c9f", X"9c97", 
X"9c8f", X"9c87", X"9c7f", X"9c77", X"9c6f", X"9c67", X"9c60", X"9c58", 
X"9c50", X"9c48", X"9c40", X"9c38", X"9c30", X"9c28", X"9c21", X"9c19", 
X"9c11", X"9c09", X"9c01", X"9bf9", X"9bf1", X"9bea", X"9be2", X"9bda", 
X"9bd2", X"9bca", X"9bc2", X"9bbb", X"9bb3", X"9bab", X"9ba3", X"9b9b", 
X"9b94", X"9b8c", X"9b84", X"9b7c", X"9b75", X"9b6d", X"9b65", X"9b5d", 
X"9b55", X"9b4e", X"9b46", X"9b3e", X"9b36", X"9b2f", X"9b27", X"9b1f", 
X"9b17", X"9b10", X"9b08", X"9b00", X"9af9", X"9af1", X"9ae9", X"9ae1", 
X"9ada", X"9ad2", X"9aca", X"9ac3", X"9abb", X"9ab3", X"9aac", X"9aa4", 
X"9a9c", X"9a95", X"9a8d", X"9a85", X"9a7e", X"9a76", X"9a6e", X"9a67", 
X"9a5f", X"9a57", X"9a50", X"9a48", X"9a40", X"9a39", X"9a31", X"9a2a", 
X"9a22", X"9a1a", X"9a13", X"9a0b", X"9a04", X"99fc", X"99f4", X"99ed", 
X"99e5", X"99de", X"99d6", X"99cf", X"99c7", X"99bf", X"99b8", X"99b0", 
X"99a9", X"99a1", X"999a", X"9992", X"998b", X"9983", X"997c", X"9974", 
X"996d", X"9965", X"995d", X"9956", X"994e", X"9947", X"993f", X"9938", 
X"9930", X"9929", X"9922", X"991a", X"9913", X"990b", X"9904", X"98fc", 
X"98f5", X"98ed", X"98e6", X"98de", X"98d7", X"98d0", X"98c8", X"98c1", 
X"98b9", X"98b2", X"98aa", X"98a3", X"989c", X"9894", X"988d", X"9885", 
X"987e", X"9877", X"986f", X"9868", X"9860", X"9859", X"9852", X"984a", 
X"9843", X"983c", X"9834", X"982d", X"9826", X"981e", X"9817", X"9810", 
X"9808", X"9801", X"97fa", X"97f2", X"97eb", X"97e4", X"97dc", X"97d5", 
X"97ce", X"97c6", X"97bf", X"97b8", X"97b0", X"97a9", X"97a2", X"979b", 
X"9793", X"978c", X"9785", X"977e", X"9776", X"976f", X"9768", X"9761", 
X"9759", X"9752", X"974b", X"9744", X"973c", X"9735", X"972e", X"9727", 
X"9720", X"9718", X"9711", X"970a", X"9703", X"96fc", X"96f4", X"96ed", 
X"96e6", X"96df", X"96d8", X"96d1", X"96c9", X"96c2", X"96bb", X"96b4", 
X"96ad", X"96a6", X"969f", X"9697", X"9690", X"9689", X"9682", X"967b", 
X"9674", X"966d", X"9666", X"965f", X"9657", X"9650", X"9649", X"9642", 
X"963b", X"9634", X"962d", X"9626", X"961f", X"9618", X"9611", X"960a", 
X"9603", X"95fc", X"95f5", X"95ee", X"95e6", X"95df", X"95d8", X"95d1", 
X"95ca", X"95c3", X"95bc", X"95b5", X"95ae", X"95a7", X"95a0", X"9599", 
X"9592", X"958b", X"9584", X"957d", X"9577", X"9570", X"9569", X"9562", 
X"955b", X"9554", X"954d", X"9546", X"953f", X"9538", X"9531", X"952a", 
X"9523", X"951c", X"9515", X"950e", X"9508", X"9501", X"94fa", X"94f3", 
X"94ec", X"94e5", X"94de", X"94d7", X"94d0", X"94ca", X"94c3", X"94bc", 
X"94b5", X"94ae", X"94a7", X"94a1", X"949a", X"9493", X"948c", X"9485", 
X"947e", X"9478", X"9471", X"946a", X"9463", X"945c", X"9456", X"944f", 
X"9448", X"9441", X"943a", X"9434", X"942d", X"9426", X"941f", X"9419", 
X"9412", X"940b", X"9404", X"93fe", X"93f7", X"93f0", X"93e9", X"93e3", 
X"93dc", X"93d5", X"93ce", X"93c8", X"93c1", X"93ba", X"93b4", X"93ad", 
X"93a6", X"939f", X"9399", X"9392", X"938b", X"9385", X"937e", X"9377", 
X"9371", X"936a", X"9363", X"935d", X"9356", X"9350", X"9349", X"9342", 
X"933c", X"9335", X"932e", X"9328", X"9321", X"931b", X"9314", X"930d", 
X"9307", X"9300", X"92fa", X"92f3", X"92ec", X"92e6", X"92df", X"92d9", 
X"92d2", X"92cc", X"92c5", X"92bf", X"92b8", X"92b1", X"92ab", X"92a4", 
X"929e", X"9297", X"9291", X"928a", X"9284", X"927d", X"9277", X"9270", 
X"926a", X"9263", X"925d", X"9256", X"9250", X"9249", X"9243", X"923c", 
X"9236", X"922f", X"9229", X"9223", X"921c", X"9216", X"920f", X"9209", 
X"9202", X"91fc", X"91f6", X"91ef", X"91e9", X"91e2", X"91dc", X"91d6", 
X"91cf", X"91c9", X"91c2", X"91bc", X"91b6", X"91af", X"91a9", X"91a2", 
X"919c", X"9196", X"918f", X"9189", X"9183", X"917c", X"9176", X"9170", 
X"9169", X"9163", X"915d", X"9156", X"9150", X"914a", X"9143", X"913d", 
X"9137", X"9131", X"912a", X"9124", X"911e", X"9117", X"9111", X"910b", 
X"9105", X"90fe", X"90f8", X"90f2", X"90ec", X"90e5", X"90df", X"90d9", 
X"90d3", X"90cc", X"90c6", X"90c0", X"90ba", X"90b4", X"90ad", X"90a7", 
X"90a1", X"909b", X"9095", X"908e", X"9088", X"9082", X"907c", X"9076", 
X"9070", X"9069", X"9063", X"905d", X"9057", X"9051", X"904b", X"9045", 
X"903e", X"9038", X"9032", X"902c", X"9026", X"9020", X"901a", X"9014", 
X"900e", X"9007", X"9001", X"8ffb", X"8ff5", X"8fef", X"8fe9", X"8fe3", 
X"8fdd", X"8fd7", X"8fd1", X"8fcb", X"8fc5", X"8fbf", X"8fb9", X"8fb3", 
X"8fad", X"8fa7", X"8fa1", X"8f9b", X"8f95", X"8f8f", X"8f89", X"8f83", 
X"8f7d", X"8f77", X"8f71", X"8f6b", X"8f65", X"8f5f", X"8f59", X"8f53", 
X"8f4d", X"8f47", X"8f41", X"8f3b", X"8f35", X"8f2f", X"8f29", X"8f23", 
X"8f1d", X"8f17", X"8f11", X"8f0b", X"8f06", X"8f00", X"8efa", X"8ef4", 
X"8eee", X"8ee8", X"8ee2", X"8edc", X"8ed6", X"8ed1", X"8ecb", X"8ec5", 
X"8ebf", X"8eb9", X"8eb3", X"8ead", X"8ea8", X"8ea2", X"8e9c", X"8e96", 
X"8e90", X"8e8a", X"8e85", X"8e7f", X"8e79", X"8e73", X"8e6d", X"8e68", 
X"8e62", X"8e5c", X"8e56", X"8e50", X"8e4b", X"8e45", X"8e3f", X"8e39", 
X"8e34", X"8e2e", X"8e28", X"8e22", X"8e1d", X"8e17", X"8e11", X"8e0b", 
X"8e06", X"8e00", X"8dfa", X"8df5", X"8def", X"8de9", X"8de4", X"8dde", 
X"8dd8", X"8dd2", X"8dcd", X"8dc7", X"8dc1", X"8dbc", X"8db6", X"8db0", 
X"8dab", X"8da5", X"8da0", X"8d9a", X"8d94", X"8d8f", X"8d89", X"8d83", 
X"8d7e", X"8d78", X"8d73", X"8d6d", X"8d67", X"8d62", X"8d5c", X"8d57", 
X"8d51", X"8d4b", X"8d46", X"8d40", X"8d3b", X"8d35", X"8d30", X"8d2a", 
X"8d24", X"8d1f", X"8d19", X"8d14", X"8d0e", X"8d09", X"8d03", X"8cfe", 
X"8cf8", X"8cf3", X"8ced", X"8ce8", X"8ce2", X"8cdd", X"8cd7", X"8cd2", 
X"8ccc", X"8cc7", X"8cc1", X"8cbc", X"8cb6", X"8cb1", X"8cab", X"8ca6", 
X"8ca1", X"8c9b", X"8c96", X"8c90", X"8c8b", X"8c85", X"8c80", X"8c7b", 
X"8c75", X"8c70", X"8c6a", X"8c65", X"8c60", X"8c5a", X"8c55", X"8c4f", 
X"8c4a", X"8c45", X"8c3f", X"8c3a", X"8c35", X"8c2f", X"8c2a", X"8c25", 
X"8c1f", X"8c1a", X"8c15", X"8c0f", X"8c0a", X"8c05", X"8bff", X"8bfa", 
X"8bf5", X"8bef", X"8bea", X"8be5", X"8bdf", X"8bda", X"8bd5", X"8bd0", 
X"8bca", X"8bc5", X"8bc0", X"8bbb", X"8bb5", X"8bb0", X"8bab", X"8ba6", 
X"8ba0", X"8b9b", X"8b96", X"8b91", X"8b8b", X"8b86", X"8b81", X"8b7c", 
X"8b77", X"8b71", X"8b6c", X"8b67", X"8b62", X"8b5d", X"8b58", X"8b52", 
X"8b4d", X"8b48", X"8b43", X"8b3e", X"8b39", X"8b33", X"8b2e", X"8b29", 
X"8b24", X"8b1f", X"8b1a", X"8b15", X"8b10", X"8b0a", X"8b05", X"8b00", 
X"8afb", X"8af6", X"8af1", X"8aec", X"8ae7", X"8ae2", X"8add", X"8ad8", 
X"8ad3", X"8ace", X"8ac8", X"8ac3", X"8abe", X"8ab9", X"8ab4", X"8aaf", 
X"8aaa", X"8aa5", X"8aa0", X"8a9b", X"8a96", X"8a91", X"8a8c", X"8a87", 
X"8a82", X"8a7d", X"8a78", X"8a73", X"8a6e", X"8a69", X"8a64", X"8a5f", 
X"8a5a", X"8a56", X"8a51", X"8a4c", X"8a47", X"8a42", X"8a3d", X"8a38", 
X"8a33", X"8a2e", X"8a29", X"8a24", X"8a1f", X"8a1a", X"8a16", X"8a11", 
X"8a0c", X"8a07", X"8a02", X"89fd", X"89f8", X"89f3", X"89ef", X"89ea", 
X"89e5", X"89e0", X"89db", X"89d6", X"89d2", X"89cd", X"89c8", X"89c3", 
X"89be", X"89ba", X"89b5", X"89b0", X"89ab", X"89a6", X"89a2", X"899d", 
X"8998", X"8993", X"898e", X"898a", X"8985", X"8980", X"897b", X"8977", 
X"8972", X"896d", X"8968", X"8964", X"895f", X"895a", X"8956", X"8951", 
X"894c", X"8947", X"8943", X"893e", X"8939", X"8935", X"8930", X"892b", 
X"8927", X"8922", X"891d", X"8919", X"8914", X"890f", X"890b", X"8906", 
X"8902", X"88fd", X"88f8", X"88f4", X"88ef", X"88ea", X"88e6", X"88e1", 
X"88dd", X"88d8", X"88d3", X"88cf", X"88ca", X"88c6", X"88c1", X"88bd", 
X"88b8", X"88b3", X"88af", X"88aa", X"88a6", X"88a1", X"889d", X"8898", 
X"8894", X"888f", X"888b", X"8886", X"8882", X"887d", X"8879", X"8874", 
X"8870", X"886b", X"8867", X"8862", X"885e", X"8859", X"8855", X"8850", 
X"884c", X"8847", X"8843", X"883f", X"883a", X"8836", X"8831", X"882d", 
X"8828", X"8824", X"8820", X"881b", X"8817", X"8812", X"880e", X"880a", 
X"8805", X"8801", X"87fd", X"87f8", X"87f4", X"87ef", X"87eb", X"87e7", 
X"87e2", X"87de", X"87da", X"87d5", X"87d1", X"87cd", X"87c8", X"87c4", 
X"87c0", X"87bb", X"87b7", X"87b3", X"87af", X"87aa", X"87a6", X"87a2", 
X"879d", X"8799", X"8795", X"8791", X"878c", X"8788", X"8784", X"8780", 
X"877b", X"8777", X"8773", X"876f", X"876b", X"8766", X"8762", X"875e", 
X"875a", X"8756", X"8751", X"874d", X"8749", X"8745", X"8741", X"873c", 
X"8738", X"8734", X"8730", X"872c", X"8728", X"8724", X"871f", X"871b", 
X"8717", X"8713", X"870f", X"870b", X"8707", X"8703", X"86ff", X"86fa", 
X"86f6", X"86f2", X"86ee", X"86ea", X"86e6", X"86e2", X"86de", X"86da", 
X"86d6", X"86d2", X"86ce", X"86ca", X"86c6", X"86c2", X"86be", X"86ba", 
X"86b6", X"86b2", X"86ad", X"86a9", X"86a5", X"86a1", X"869e", X"869a", 
X"8696", X"8692", X"868e", X"868a", X"8686", X"8682", X"867e", X"867a", 
X"8676", X"8672", X"866e", X"866a", X"8666", X"8662", X"865e", X"865a", 
X"8656", X"8653", X"864f", X"864b", X"8647", X"8643", X"863f", X"863b", 
X"8637", X"8634", X"8630", X"862c", X"8628", X"8624", X"8620", X"861c", 
X"8619", X"8615", X"8611", X"860d", X"8609", X"8605", X"8602", X"85fe", 
X"85fa", X"85f6", X"85f2", X"85ef", X"85eb", X"85e7", X"85e3", X"85e0", 
X"85dc", X"85d8", X"85d4", X"85d1", X"85cd", X"85c9", X"85c5", X"85c2", 
X"85be", X"85ba", X"85b7", X"85b3", X"85af", X"85ab", X"85a8", X"85a4", 
X"85a0", X"859d", X"8599", X"8595", X"8592", X"858e", X"858a", X"8587", 
X"8583", X"857f", X"857c", X"8578", X"8574", X"8571", X"856d", X"856a", 
X"8566", X"8562", X"855f", X"855b", X"8558", X"8554", X"8550", X"854d", 
X"8549", X"8546", X"8542", X"853f", X"853b", X"8537", X"8534", X"8530", 
X"852d", X"8529", X"8526", X"8522", X"851f", X"851b", X"8518", X"8514", 
X"8511", X"850d", X"850a", X"8506", X"8503", X"84ff", X"84fc", X"84f8", 
X"84f5", X"84f1", X"84ee", X"84ea", X"84e7", X"84e4", X"84e0", X"84dd", 
X"84d9", X"84d6", X"84d2", X"84cf", X"84cc", X"84c8", X"84c5", X"84c1", 
X"84be", X"84bb", X"84b7", X"84b4", X"84b0", X"84ad", X"84aa", X"84a6", 
X"84a3", X"84a0", X"849c", X"8499", X"8496", X"8492", X"848f", X"848c", 
X"8488", X"8485", X"8482", X"847e", X"847b", X"8478", X"8475", X"8471", 
X"846e", X"846b", X"8467", X"8464", X"8461", X"845e", X"845a", X"8457", 
X"8454", X"8451", X"844d", X"844a", X"8447", X"8444", X"8441", X"843d", 
X"843a", X"8437", X"8434", X"8431", X"842d", X"842a", X"8427", X"8424", 
X"8421", X"841d", X"841a", X"8417", X"8414", X"8411", X"840e", X"840b", 
X"8407", X"8404", X"8401", X"83fe", X"83fb", X"83f8", X"83f5", X"83f2", 
X"83ef", X"83ec", X"83e8", X"83e5", X"83e2", X"83df", X"83dc", X"83d9", 
X"83d6", X"83d3", X"83d0", X"83cd", X"83ca", X"83c7", X"83c4", X"83c1", 
X"83be", X"83bb", X"83b8", X"83b5", X"83b2", X"83af", X"83ac", X"83a9", 
X"83a6", X"83a3", X"83a0", X"839d", X"839a", X"8397", X"8394", X"8391", 
X"838e", X"838b", X"8388", X"8385", X"8382", X"837f", X"837d", X"837a", 
X"8377", X"8374", X"8371", X"836e", X"836b", X"8368", X"8365", X"8362", 
X"8360", X"835d", X"835a", X"8357", X"8354", X"8351", X"834f", X"834c", 
X"8349", X"8346", X"8343", X"8340", X"833e", X"833b", X"8338", X"8335", 
X"8332", X"8330", X"832d", X"832a", X"8327", X"8324", X"8322", X"831f", 
X"831c", X"8319", X"8317", X"8314", X"8311", X"830e", X"830c", X"8309", 
X"8306", X"8304", X"8301", X"82fe", X"82fb", X"82f9", X"82f6", X"82f3", 
X"82f1", X"82ee", X"82eb", X"82e9", X"82e6", X"82e3", X"82e1", X"82de", 
X"82db", X"82d9", X"82d6", X"82d4", X"82d1", X"82ce", X"82cc", X"82c9", 
X"82c6", X"82c4", X"82c1", X"82bf", X"82bc", X"82ba", X"82b7", X"82b4", 
X"82b2", X"82af", X"82ad", X"82aa", X"82a8", X"82a5", X"82a3", X"82a0", 
X"829d", X"829b", X"8298", X"8296", X"8293", X"8291", X"828e", X"828c", 
X"8289", X"8287", X"8284", X"8282", X"827f", X"827d", X"827b", X"8278", 
X"8276", X"8273", X"8271", X"826e", X"826c", X"8269", X"8267", X"8265", 
X"8262", X"8260", X"825d", X"825b", X"8259", X"8256", X"8254", X"8251", 
X"824f", X"824d", X"824a", X"8248", X"8246", X"8243", X"8241", X"823e", 
X"823c", X"823a", X"8237", X"8235", X"8233", X"8231", X"822e", X"822c", 
X"822a", X"8227", X"8225", X"8223", X"8220", X"821e", X"821c", X"821a", 
X"8217", X"8215", X"8213", X"8211", X"820e", X"820c", X"820a", X"8208", 
X"8205", X"8203", X"8201", X"81ff", X"81fd", X"81fa", X"81f8", X"81f6", 
X"81f4", X"81f2", X"81ef", X"81ed", X"81eb", X"81e9", X"81e7", X"81e5", 
X"81e2", X"81e0", X"81de", X"81dc", X"81da", X"81d8", X"81d6", X"81d3", 
X"81d1", X"81cf", X"81cd", X"81cb", X"81c9", X"81c7", X"81c5", X"81c3", 
X"81c1", X"81bf", X"81bd", X"81ba", X"81b8", X"81b6", X"81b4", X"81b2", 
X"81b0", X"81ae", X"81ac", X"81aa", X"81a8", X"81a6", X"81a4", X"81a2", 
X"81a0", X"819e", X"819c", X"819a", X"8198", X"8196", X"8194", X"8192", 
X"8190", X"818e", X"818c", X"818a", X"8188", X"8187", X"8185", X"8183", 
X"8181", X"817f", X"817d", X"817b", X"8179", X"8177", X"8175", X"8173", 
X"8172", X"8170", X"816e", X"816c", X"816a", X"8168", X"8166", X"8165", 
X"8163", X"8161", X"815f", X"815d", X"815b", X"815a", X"8158", X"8156", 
X"8154", X"8152", X"8150", X"814f", X"814d", X"814b", X"8149", X"8148", 
X"8146", X"8144", X"8142", X"8140", X"813f", X"813d", X"813b", X"813a", 
X"8138", X"8136", X"8134", X"8133", X"8131", X"812f", X"812d", X"812c", 
X"812a", X"8128", X"8127", X"8125", X"8123", X"8122", X"8120", X"811e", 
X"811d", X"811b", X"8119", X"8118", X"8116", X"8115", X"8113", X"8111", 
X"8110", X"810e", X"810c", X"810b", X"8109", X"8108", X"8106", X"8104", 
X"8103", X"8101", X"8100", X"80fe", X"80fd", X"80fb", X"80fa", X"80f8", 
X"80f6", X"80f5", X"80f3", X"80f2", X"80f0", X"80ef", X"80ed", X"80ec", 
X"80ea", X"80e9", X"80e7", X"80e6", X"80e4", X"80e3", X"80e1", X"80e0", 
X"80de", X"80dd", X"80dc", X"80da", X"80d9", X"80d7", X"80d6", X"80d4", 
X"80d3", X"80d1", X"80d0", X"80cf", X"80cd", X"80cc", X"80ca", X"80c9", 
X"80c8", X"80c6", X"80c5", X"80c4", X"80c2", X"80c1", X"80bf", X"80be", 
X"80bd", X"80bb", X"80ba", X"80b9", X"80b7", X"80b6", X"80b5", X"80b3", 
X"80b2", X"80b1", X"80b0", X"80ae", X"80ad", X"80ac", X"80aa", X"80a9", 
X"80a8", X"80a7", X"80a5", X"80a4", X"80a3", X"80a2", X"80a0", X"809f", 
X"809e", X"809d", X"809b", X"809a", X"8099", X"8098", X"8096", X"8095", 
X"8094", X"8093", X"8092", X"8091", X"808f", X"808e", X"808d", X"808c", 
X"808b", X"808a", X"8088", X"8087", X"8086", X"8085", X"8084", X"8083", 
X"8082", X"8080", X"807f", X"807e", X"807d", X"807c", X"807b", X"807a", 
X"8079", X"8078", X"8077", X"8076", X"8075", X"8073", X"8072", X"8071", 
X"8070", X"806f", X"806e", X"806d", X"806c", X"806b", X"806a", X"8069", 
X"8068", X"8067", X"8066", X"8065", X"8064", X"8063", X"8062", X"8061", 
X"8060", X"805f", X"805e", X"805d", X"805d", X"805c", X"805b", X"805a", 
X"8059", X"8058", X"8057", X"8056", X"8055", X"8054", X"8053", X"8052", 
X"8052", X"8051", X"8050", X"804f", X"804e", X"804d", X"804c", X"804b", 
X"804b", X"804a", X"8049", X"8048", X"8047", X"8046", X"8046", X"8045", 
X"8044", X"8043", X"8042", X"8042", X"8041", X"8040", X"803f", X"803e", 
X"803e", X"803d", X"803c", X"803b", X"803b", X"803a", X"8039", X"8038", 
X"8038", X"8037", X"8036", X"8035", X"8035", X"8034", X"8033", X"8033", 
X"8032", X"8031", X"8031", X"8030", X"802f", X"802f", X"802e", X"802d", 
X"802d", X"802c", X"802b", X"802b", X"802a", X"8029", X"8029", X"8028", 
X"8027", X"8027", X"8026", X"8026", X"8025", X"8024", X"8024", X"8023", 
X"8023", X"8022", X"8022", X"8021", X"8020", X"8020", X"801f", X"801f", 
X"801e", X"801e", X"801d", X"801d", X"801c", X"801c", X"801b", X"801b", 
X"801a", X"801a", X"8019", X"8019", X"8018", X"8018", X"8017", X"8017", 
X"8016", X"8016", X"8015", X"8015", X"8014", X"8014", X"8014", X"8013", 
X"8013", X"8012", X"8012", X"8011", X"8011", X"8011", X"8010", X"8010", 
X"800f", X"800f", X"800f", X"800e", X"800e", X"800e", X"800d", X"800d", 
X"800c", X"800c", X"800c", X"800b", X"800b", X"800b", X"800a", X"800a", 
X"800a", X"800a", X"8009", X"8009", X"8009", X"8008", X"8008", X"8008", 
X"8008", X"8007", X"8007", X"8007", X"8007", X"8006", X"8006", X"8006", 
X"8006", X"8005", X"8005", X"8005", X"8005", X"8004", X"8004", X"8004", 
X"8004", X"8004", X"8003", X"8003", X"8003", X"8003", X"8003", X"8003", 
X"8002", X"8002", X"8002", X"8002", X"8002", X"8002", X"8002", X"8002", 
X"8001", X"8001", X"8001", X"8001", X"8001", X"8001", X"8001", X"8001", 
X"8001", X"8001", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8001", 
X"8001", X"8001", X"8001", X"8001", X"8001", X"8001", X"8001", X"8001", 
X"8001", X"8002", X"8002", X"8002", X"8002", X"8002", X"8002", X"8002", 
X"8002", X"8003", X"8003", X"8003", X"8003", X"8003", X"8003", X"8004", 
X"8004", X"8004", X"8004", X"8004", X"8005", X"8005", X"8005", X"8005", 
X"8006", X"8006", X"8006", X"8006", X"8007", X"8007", X"8007", X"8007", 
X"8008", X"8008", X"8008", X"8008", X"8009", X"8009", X"8009", X"800a", 
X"800a", X"800a", X"800a", X"800b", X"800b", X"800b", X"800c", X"800c", 
X"800c", X"800d", X"800d", X"800e", X"800e", X"800e", X"800f", X"800f", 
X"800f", X"8010", X"8010", X"8011", X"8011", X"8011", X"8012", X"8012", 
X"8013", X"8013", X"8014", X"8014", X"8014", X"8015", X"8015", X"8016", 
X"8016", X"8017", X"8017", X"8018", X"8018", X"8019", X"8019", X"801a", 
X"801a", X"801b", X"801b", X"801c", X"801c", X"801d", X"801d", X"801e", 
X"801e", X"801f", X"801f", X"8020", X"8020", X"8021", X"8022", X"8022", 
X"8023", X"8023", X"8024", X"8024", X"8025", X"8026", X"8026", X"8027", 
X"8027", X"8028", X"8029", X"8029", X"802a", X"802b", X"802b", X"802c", 
X"802d", X"802d", X"802e", X"802f", X"802f", X"8030", X"8031", X"8031", 
X"8032", X"8033", X"8033", X"8034", X"8035", X"8035", X"8036", X"8037", 
X"8038", X"8038", X"8039", X"803a", X"803b", X"803b", X"803c", X"803d", 
X"803e", X"803e", X"803f", X"8040", X"8041", X"8042", X"8042", X"8043", 
X"8044", X"8045", X"8046", X"8046", X"8047", X"8048", X"8049", X"804a", 
X"804b", X"804b", X"804c", X"804d", X"804e", X"804f", X"8050", X"8051", 
X"8052", X"8052", X"8053", X"8054", X"8055", X"8056", X"8057", X"8058", 
X"8059", X"805a", X"805b", X"805c", X"805d", X"805d", X"805e", X"805f", 
X"8060", X"8061", X"8062", X"8063", X"8064", X"8065", X"8066", X"8067", 
X"8068", X"8069", X"806a", X"806b", X"806c", X"806d", X"806e", X"806f", 
X"8070", X"8071", X"8072", X"8073", X"8075", X"8076", X"8077", X"8078", 
X"8079", X"807a", X"807b", X"807c", X"807d", X"807e", X"807f", X"8080", 
X"8082", X"8083", X"8084", X"8085", X"8086", X"8087", X"8088", X"808a", 
X"808b", X"808c", X"808d", X"808e", X"808f", X"8091", X"8092", X"8093", 
X"8094", X"8095", X"8096", X"8098", X"8099", X"809a", X"809b", X"809d", 
X"809e", X"809f", X"80a0", X"80a2", X"80a3", X"80a4", X"80a5", X"80a7", 
X"80a8", X"80a9", X"80aa", X"80ac", X"80ad", X"80ae", X"80b0", X"80b1", 
X"80b2", X"80b3", X"80b5", X"80b6", X"80b7", X"80b9", X"80ba", X"80bb", 
X"80bd", X"80be", X"80bf", X"80c1", X"80c2", X"80c4", X"80c5", X"80c6", 
X"80c8", X"80c9", X"80ca", X"80cc", X"80cd", X"80cf", X"80d0", X"80d1", 
X"80d3", X"80d4", X"80d6", X"80d7", X"80d9", X"80da", X"80dc", X"80dd", 
X"80de", X"80e0", X"80e1", X"80e3", X"80e4", X"80e6", X"80e7", X"80e9", 
X"80ea", X"80ec", X"80ed", X"80ef", X"80f0", X"80f2", X"80f3", X"80f5", 
X"80f6", X"80f8", X"80fa", X"80fb", X"80fd", X"80fe", X"8100", X"8101", 
X"8103", X"8104", X"8106", X"8108", X"8109", X"810b", X"810c", X"810e", 
X"8110", X"8111", X"8113", X"8115", X"8116", X"8118", X"8119", X"811b", 
X"811d", X"811e", X"8120", X"8122", X"8123", X"8125", X"8127", X"8128", 
X"812a", X"812c", X"812d", X"812f", X"8131", X"8133", X"8134", X"8136", 
X"8138", X"813a", X"813b", X"813d", X"813f", X"8140", X"8142", X"8144", 
X"8146", X"8148", X"8149", X"814b", X"814d", X"814f", X"8150", X"8152", 
X"8154", X"8156", X"8158", X"815a", X"815b", X"815d", X"815f", X"8161", 
X"8163", X"8165", X"8166", X"8168", X"816a", X"816c", X"816e", X"8170", 
X"8172", X"8173", X"8175", X"8177", X"8179", X"817b", X"817d", X"817f", 
X"8181", X"8183", X"8185", X"8187", X"8188", X"818a", X"818c", X"818e", 
X"8190", X"8192", X"8194", X"8196", X"8198", X"819a", X"819c", X"819e", 
X"81a0", X"81a2", X"81a4", X"81a6", X"81a8", X"81aa", X"81ac", X"81ae", 
X"81b0", X"81b2", X"81b4", X"81b6", X"81b8", X"81ba", X"81bd", X"81bf", 
X"81c1", X"81c3", X"81c5", X"81c7", X"81c9", X"81cb", X"81cd", X"81cf", 
X"81d1", X"81d3", X"81d6", X"81d8", X"81da", X"81dc", X"81de", X"81e0", 
X"81e2", X"81e5", X"81e7", X"81e9", X"81eb", X"81ed", X"81ef", X"81f2", 
X"81f4", X"81f6", X"81f8", X"81fa", X"81fd", X"81ff", X"8201", X"8203", 
X"8205", X"8208", X"820a", X"820c", X"820e", X"8211", X"8213", X"8215", 
X"8217", X"821a", X"821c", X"821e", X"8220", X"8223", X"8225", X"8227", 
X"822a", X"822c", X"822e", X"8231", X"8233", X"8235", X"8237", X"823a", 
X"823c", X"823e", X"8241", X"8243", X"8246", X"8248", X"824a", X"824d", 
X"824f", X"8251", X"8254", X"8256", X"8259", X"825b", X"825d", X"8260", 
X"8262", X"8265", X"8267", X"8269", X"826c", X"826e", X"8271", X"8273", 
X"8276", X"8278", X"827b", X"827d", X"827f", X"8282", X"8284", X"8287", 
X"8289", X"828c", X"828e", X"8291", X"8293", X"8296", X"8298", X"829b", 
X"829d", X"82a0", X"82a3", X"82a5", X"82a8", X"82aa", X"82ad", X"82af", 
X"82b2", X"82b4", X"82b7", X"82ba", X"82bc", X"82bf", X"82c1", X"82c4", 
X"82c6", X"82c9", X"82cc", X"82ce", X"82d1", X"82d4", X"82d6", X"82d9", 
X"82db", X"82de", X"82e1", X"82e3", X"82e6", X"82e9", X"82eb", X"82ee", 
X"82f1", X"82f3", X"82f6", X"82f9", X"82fb", X"82fe", X"8301", X"8304", 
X"8306", X"8309", X"830c", X"830e", X"8311", X"8314", X"8317", X"8319", 
X"831c", X"831f", X"8322", X"8324", X"8327", X"832a", X"832d", X"8330", 
X"8332", X"8335", X"8338", X"833b", X"833e", X"8340", X"8343", X"8346", 
X"8349", X"834c", X"834f", X"8351", X"8354", X"8357", X"835a", X"835d", 
X"8360", X"8362", X"8365", X"8368", X"836b", X"836e", X"8371", X"8374", 
X"8377", X"837a", X"837d", X"837f", X"8382", X"8385", X"8388", X"838b", 
X"838e", X"8391", X"8394", X"8397", X"839a", X"839d", X"83a0", X"83a3", 
X"83a6", X"83a9", X"83ac", X"83af", X"83b2", X"83b5", X"83b8", X"83bb", 
X"83be", X"83c1", X"83c4", X"83c7", X"83ca", X"83cd", X"83d0", X"83d3", 
X"83d6", X"83d9", X"83dc", X"83df", X"83e2", X"83e5", X"83e8", X"83ec", 
X"83ef", X"83f2", X"83f5", X"83f8", X"83fb", X"83fe", X"8401", X"8404", 
X"8407", X"840b", X"840e", X"8411", X"8414", X"8417", X"841a", X"841d", 
X"8421", X"8424", X"8427", X"842a", X"842d", X"8431", X"8434", X"8437", 
X"843a", X"843d", X"8441", X"8444", X"8447", X"844a", X"844d", X"8451", 
X"8454", X"8457", X"845a", X"845e", X"8461", X"8464", X"8467", X"846b", 
X"846e", X"8471", X"8475", X"8478", X"847b", X"847e", X"8482", X"8485", 
X"8488", X"848c", X"848f", X"8492", X"8496", X"8499", X"849c", X"84a0", 
X"84a3", X"84a6", X"84aa", X"84ad", X"84b0", X"84b4", X"84b7", X"84bb", 
X"84be", X"84c1", X"84c5", X"84c8", X"84cc", X"84cf", X"84d2", X"84d6", 
X"84d9", X"84dd", X"84e0", X"84e4", X"84e7", X"84ea", X"84ee", X"84f1", 
X"84f5", X"84f8", X"84fc", X"84ff", X"8503", X"8506", X"850a", X"850d", 
X"8511", X"8514", X"8518", X"851b", X"851f", X"8522", X"8526", X"8529", 
X"852d", X"8530", X"8534", X"8537", X"853b", X"853f", X"8542", X"8546", 
X"8549", X"854d", X"8550", X"8554", X"8558", X"855b", X"855f", X"8562", 
X"8566", X"856a", X"856d", X"8571", X"8574", X"8578", X"857c", X"857f", 
X"8583", X"8587", X"858a", X"858e", X"8592", X"8595", X"8599", X"859d", 
X"85a0", X"85a4", X"85a8", X"85ab", X"85af", X"85b3", X"85b7", X"85ba", 
X"85be", X"85c2", X"85c5", X"85c9", X"85cd", X"85d1", X"85d4", X"85d8", 
X"85dc", X"85e0", X"85e3", X"85e7", X"85eb", X"85ef", X"85f2", X"85f6", 
X"85fa", X"85fe", X"8602", X"8605", X"8609", X"860d", X"8611", X"8615", 
X"8619", X"861c", X"8620", X"8624", X"8628", X"862c", X"8630", X"8634", 
X"8637", X"863b", X"863f", X"8643", X"8647", X"864b", X"864f", X"8653", 
X"8656", X"865a", X"865e", X"8662", X"8666", X"866a", X"866e", X"8672", 
X"8676", X"867a", X"867e", X"8682", X"8686", X"868a", X"868e", X"8692", 
X"8696", X"869a", X"869e", X"86a1", X"86a5", X"86a9", X"86ad", X"86b2", 
X"86b6", X"86ba", X"86be", X"86c2", X"86c6", X"86ca", X"86ce", X"86d2", 
X"86d6", X"86da", X"86de", X"86e2", X"86e6", X"86ea", X"86ee", X"86f2", 
X"86f6", X"86fa", X"86ff", X"8703", X"8707", X"870b", X"870f", X"8713", 
X"8717", X"871b", X"871f", X"8724", X"8728", X"872c", X"8730", X"8734", 
X"8738", X"873c", X"8741", X"8745", X"8749", X"874d", X"8751", X"8756", 
X"875a", X"875e", X"8762", X"8766", X"876b", X"876f", X"8773", X"8777", 
X"877b", X"8780", X"8784", X"8788", X"878c", X"8791", X"8795", X"8799", 
X"879d", X"87a2", X"87a6", X"87aa", X"87af", X"87b3", X"87b7", X"87bb", 
X"87c0", X"87c4", X"87c8", X"87cd", X"87d1", X"87d5", X"87da", X"87de", 
X"87e2", X"87e7", X"87eb", X"87ef", X"87f4", X"87f8", X"87fd", X"8801", 
X"8805", X"880a", X"880e", X"8812", X"8817", X"881b", X"8820", X"8824", 
X"8828", X"882d", X"8831", X"8836", X"883a", X"883f", X"8843", X"8847", 
X"884c", X"8850", X"8855", X"8859", X"885e", X"8862", X"8867", X"886b", 
X"8870", X"8874", X"8879", X"887d", X"8882", X"8886", X"888b", X"888f", 
X"8894", X"8898", X"889d", X"88a1", X"88a6", X"88aa", X"88af", X"88b3", 
X"88b8", X"88bd", X"88c1", X"88c6", X"88ca", X"88cf", X"88d3", X"88d8", 
X"88dd", X"88e1", X"88e6", X"88ea", X"88ef", X"88f4", X"88f8", X"88fd", 
X"8902", X"8906", X"890b", X"890f", X"8914", X"8919", X"891d", X"8922", 
X"8927", X"892b", X"8930", X"8935", X"8939", X"893e", X"8943", X"8947", 
X"894c", X"8951", X"8956", X"895a", X"895f", X"8964", X"8968", X"896d", 
X"8972", X"8977", X"897b", X"8980", X"8985", X"898a", X"898e", X"8993", 
X"8998", X"899d", X"89a2", X"89a6", X"89ab", X"89b0", X"89b5", X"89ba", 
X"89be", X"89c3", X"89c8", X"89cd", X"89d2", X"89d6", X"89db", X"89e0", 
X"89e5", X"89ea", X"89ef", X"89f3", X"89f8", X"89fd", X"8a02", X"8a07", 
X"8a0c", X"8a11", X"8a16", X"8a1a", X"8a1f", X"8a24", X"8a29", X"8a2e", 
X"8a33", X"8a38", X"8a3d", X"8a42", X"8a47", X"8a4c", X"8a51", X"8a56", 
X"8a5a", X"8a5f", X"8a64", X"8a69", X"8a6e", X"8a73", X"8a78", X"8a7d", 
X"8a82", X"8a87", X"8a8c", X"8a91", X"8a96", X"8a9b", X"8aa0", X"8aa5", 
X"8aaa", X"8aaf", X"8ab4", X"8ab9", X"8abe", X"8ac3", X"8ac8", X"8ace", 
X"8ad3", X"8ad8", X"8add", X"8ae2", X"8ae7", X"8aec", X"8af1", X"8af6", 
X"8afb", X"8b00", X"8b05", X"8b0a", X"8b10", X"8b15", X"8b1a", X"8b1f", 
X"8b24", X"8b29", X"8b2e", X"8b33", X"8b39", X"8b3e", X"8b43", X"8b48", 
X"8b4d", X"8b52", X"8b58", X"8b5d", X"8b62", X"8b67", X"8b6c", X"8b71", 
X"8b77", X"8b7c", X"8b81", X"8b86", X"8b8b", X"8b91", X"8b96", X"8b9b", 
X"8ba0", X"8ba6", X"8bab", X"8bb0", X"8bb5", X"8bbb", X"8bc0", X"8bc5", 
X"8bca", X"8bd0", X"8bd5", X"8bda", X"8bdf", X"8be5", X"8bea", X"8bef", 
X"8bf5", X"8bfa", X"8bff", X"8c05", X"8c0a", X"8c0f", X"8c15", X"8c1a", 
X"8c1f", X"8c25", X"8c2a", X"8c2f", X"8c35", X"8c3a", X"8c3f", X"8c45", 
X"8c4a", X"8c4f", X"8c55", X"8c5a", X"8c60", X"8c65", X"8c6a", X"8c70", 
X"8c75", X"8c7b", X"8c80", X"8c85", X"8c8b", X"8c90", X"8c96", X"8c9b", 
X"8ca1", X"8ca6", X"8cab", X"8cb1", X"8cb6", X"8cbc", X"8cc1", X"8cc7", 
X"8ccc", X"8cd2", X"8cd7", X"8cdd", X"8ce2", X"8ce8", X"8ced", X"8cf3", 
X"8cf8", X"8cfe", X"8d03", X"8d09", X"8d0e", X"8d14", X"8d19", X"8d1f", 
X"8d24", X"8d2a", X"8d30", X"8d35", X"8d3b", X"8d40", X"8d46", X"8d4b", 
X"8d51", X"8d57", X"8d5c", X"8d62", X"8d67", X"8d6d", X"8d73", X"8d78", 
X"8d7e", X"8d83", X"8d89", X"8d8f", X"8d94", X"8d9a", X"8da0", X"8da5", 
X"8dab", X"8db0", X"8db6", X"8dbc", X"8dc1", X"8dc7", X"8dcd", X"8dd2", 
X"8dd8", X"8dde", X"8de4", X"8de9", X"8def", X"8df5", X"8dfa", X"8e00", 
X"8e06", X"8e0b", X"8e11", X"8e17", X"8e1d", X"8e22", X"8e28", X"8e2e", 
X"8e34", X"8e39", X"8e3f", X"8e45", X"8e4b", X"8e50", X"8e56", X"8e5c", 
X"8e62", X"8e68", X"8e6d", X"8e73", X"8e79", X"8e7f", X"8e85", X"8e8a", 
X"8e90", X"8e96", X"8e9c", X"8ea2", X"8ea8", X"8ead", X"8eb3", X"8eb9", 
X"8ebf", X"8ec5", X"8ecb", X"8ed1", X"8ed6", X"8edc", X"8ee2", X"8ee8", 
X"8eee", X"8ef4", X"8efa", X"8f00", X"8f06", X"8f0b", X"8f11", X"8f17", 
X"8f1d", X"8f23", X"8f29", X"8f2f", X"8f35", X"8f3b", X"8f41", X"8f47", 
X"8f4d", X"8f53", X"8f59", X"8f5f", X"8f65", X"8f6b", X"8f71", X"8f77", 
X"8f7d", X"8f83", X"8f89", X"8f8f", X"8f95", X"8f9b", X"8fa1", X"8fa7", 
X"8fad", X"8fb3", X"8fb9", X"8fbf", X"8fc5", X"8fcb", X"8fd1", X"8fd7", 
X"8fdd", X"8fe3", X"8fe9", X"8fef", X"8ff5", X"8ffb", X"9001", X"9007", 
X"900e", X"9014", X"901a", X"9020", X"9026", X"902c", X"9032", X"9038", 
X"903e", X"9045", X"904b", X"9051", X"9057", X"905d", X"9063", X"9069", 
X"9070", X"9076", X"907c", X"9082", X"9088", X"908e", X"9095", X"909b", 
X"90a1", X"90a7", X"90ad", X"90b4", X"90ba", X"90c0", X"90c6", X"90cc", 
X"90d3", X"90d9", X"90df", X"90e5", X"90ec", X"90f2", X"90f8", X"90fe", 
X"9105", X"910b", X"9111", X"9117", X"911e", X"9124", X"912a", X"9131", 
X"9137", X"913d", X"9143", X"914a", X"9150", X"9156", X"915d", X"9163", 
X"9169", X"9170", X"9176", X"917c", X"9183", X"9189", X"918f", X"9196", 
X"919c", X"91a2", X"91a9", X"91af", X"91b6", X"91bc", X"91c2", X"91c9", 
X"91cf", X"91d6", X"91dc", X"91e2", X"91e9", X"91ef", X"91f6", X"91fc", 
X"9202", X"9209", X"920f", X"9216", X"921c", X"9223", X"9229", X"922f", 
X"9236", X"923c", X"9243", X"9249", X"9250", X"9256", X"925d", X"9263", 
X"926a", X"9270", X"9277", X"927d", X"9284", X"928a", X"9291", X"9297", 
X"929e", X"92a4", X"92ab", X"92b1", X"92b8", X"92bf", X"92c5", X"92cc", 
X"92d2", X"92d9", X"92df", X"92e6", X"92ec", X"92f3", X"92fa", X"9300", 
X"9307", X"930d", X"9314", X"931b", X"9321", X"9328", X"932e", X"9335", 
X"933c", X"9342", X"9349", X"9350", X"9356", X"935d", X"9363", X"936a", 
X"9371", X"9377", X"937e", X"9385", X"938b", X"9392", X"9399", X"939f", 
X"93a6", X"93ad", X"93b4", X"93ba", X"93c1", X"93c8", X"93ce", X"93d5", 
X"93dc", X"93e3", X"93e9", X"93f0", X"93f7", X"93fe", X"9404", X"940b", 
X"9412", X"9419", X"941f", X"9426", X"942d", X"9434", X"943a", X"9441", 
X"9448", X"944f", X"9456", X"945c", X"9463", X"946a", X"9471", X"9478", 
X"947e", X"9485", X"948c", X"9493", X"949a", X"94a1", X"94a7", X"94ae", 
X"94b5", X"94bc", X"94c3", X"94ca", X"94d0", X"94d7", X"94de", X"94e5", 
X"94ec", X"94f3", X"94fa", X"9501", X"9508", X"950e", X"9515", X"951c", 
X"9523", X"952a", X"9531", X"9538", X"953f", X"9546", X"954d", X"9554", 
X"955b", X"9562", X"9569", X"9570", X"9577", X"957d", X"9584", X"958b", 
X"9592", X"9599", X"95a0", X"95a7", X"95ae", X"95b5", X"95bc", X"95c3", 
X"95ca", X"95d1", X"95d8", X"95df", X"95e6", X"95ee", X"95f5", X"95fc", 
X"9603", X"960a", X"9611", X"9618", X"961f", X"9626", X"962d", X"9634", 
X"963b", X"9642", X"9649", X"9650", X"9657", X"965f", X"9666", X"966d", 
X"9674", X"967b", X"9682", X"9689", X"9690", X"9697", X"969f", X"96a6", 
X"96ad", X"96b4", X"96bb", X"96c2", X"96c9", X"96d1", X"96d8", X"96df", 
X"96e6", X"96ed", X"96f4", X"96fc", X"9703", X"970a", X"9711", X"9718", 
X"9720", X"9727", X"972e", X"9735", X"973c", X"9744", X"974b", X"9752", 
X"9759", X"9761", X"9768", X"976f", X"9776", X"977e", X"9785", X"978c", 
X"9793", X"979b", X"97a2", X"97a9", X"97b0", X"97b8", X"97bf", X"97c6", 
X"97ce", X"97d5", X"97dc", X"97e4", X"97eb", X"97f2", X"97fa", X"9801", 
X"9808", X"9810", X"9817", X"981e", X"9826", X"982d", X"9834", X"983c", 
X"9843", X"984a", X"9852", X"9859", X"9860", X"9868", X"986f", X"9877", 
X"987e", X"9885", X"988d", X"9894", X"989c", X"98a3", X"98aa", X"98b2", 
X"98b9", X"98c1", X"98c8", X"98d0", X"98d7", X"98de", X"98e6", X"98ed", 
X"98f5", X"98fc", X"9904", X"990b", X"9913", X"991a", X"9922", X"9929", 
X"9930", X"9938", X"993f", X"9947", X"994e", X"9956", X"995d", X"9965", 
X"996d", X"9974", X"997c", X"9983", X"998b", X"9992", X"999a", X"99a1", 
X"99a9", X"99b0", X"99b8", X"99bf", X"99c7", X"99cf", X"99d6", X"99de", 
X"99e5", X"99ed", X"99f4", X"99fc", X"9a04", X"9a0b", X"9a13", X"9a1a", 
X"9a22", X"9a2a", X"9a31", X"9a39", X"9a40", X"9a48", X"9a50", X"9a57", 
X"9a5f", X"9a67", X"9a6e", X"9a76", X"9a7e", X"9a85", X"9a8d", X"9a95", 
X"9a9c", X"9aa4", X"9aac", X"9ab3", X"9abb", X"9ac3", X"9aca", X"9ad2", 
X"9ada", X"9ae1", X"9ae9", X"9af1", X"9af9", X"9b00", X"9b08", X"9b10", 
X"9b17", X"9b1f", X"9b27", X"9b2f", X"9b36", X"9b3e", X"9b46", X"9b4e", 
X"9b55", X"9b5d", X"9b65", X"9b6d", X"9b75", X"9b7c", X"9b84", X"9b8c", 
X"9b94", X"9b9b", X"9ba3", X"9bab", X"9bb3", X"9bbb", X"9bc2", X"9bca", 
X"9bd2", X"9bda", X"9be2", X"9bea", X"9bf1", X"9bf9", X"9c01", X"9c09", 
X"9c11", X"9c19", X"9c21", X"9c28", X"9c30", X"9c38", X"9c40", X"9c48", 
X"9c50", X"9c58", X"9c60", X"9c67", X"9c6f", X"9c77", X"9c7f", X"9c87", 
X"9c8f", X"9c97", X"9c9f", X"9ca7", X"9caf", X"9cb7", X"9cbe", X"9cc6", 
X"9cce", X"9cd6", X"9cde", X"9ce6", X"9cee", X"9cf6", X"9cfe", X"9d06", 
X"9d0e", X"9d16", X"9d1e", X"9d26", X"9d2e", X"9d36", X"9d3e", X"9d46", 
X"9d4e", X"9d56", X"9d5e", X"9d66", X"9d6e", X"9d76", X"9d7e", X"9d86", 
X"9d8e", X"9d96", X"9d9e", X"9da6", X"9dae", X"9db6", X"9dbe", X"9dc6", 
X"9dce", X"9dd6", X"9ddf", X"9de7", X"9def", X"9df7", X"9dff", X"9e07", 
X"9e0f", X"9e17", X"9e1f", X"9e27", X"9e2f", X"9e37", X"9e40", X"9e48", 
X"9e50", X"9e58", X"9e60", X"9e68", X"9e70", X"9e78", X"9e81", X"9e89", 
X"9e91", X"9e99", X"9ea1", X"9ea9", X"9eb2", X"9eba", X"9ec2", X"9eca", 
X"9ed2", X"9eda", X"9ee3", X"9eeb", X"9ef3", X"9efb", X"9f03", X"9f0c", 
X"9f14", X"9f1c", X"9f24", X"9f2c", X"9f35", X"9f3d", X"9f45", X"9f4d", 
X"9f56", X"9f5e", X"9f66", X"9f6e", X"9f77", X"9f7f", X"9f87", X"9f8f", 
X"9f98", X"9fa0", X"9fa8", X"9fb0", X"9fb9", X"9fc1", X"9fc9", X"9fd2", 
X"9fda", X"9fe2", X"9fea", X"9ff3", X"9ffb", X"a003", X"a00c", X"a014", 
X"a01c", X"a025", X"a02d", X"a035", X"a03e", X"a046", X"a04e", X"a057", 
X"a05f", X"a067", X"a070", X"a078", X"a080", X"a089", X"a091", X"a09a", 
X"a0a2", X"a0aa", X"a0b3", X"a0bb", X"a0c4", X"a0cc", X"a0d4", X"a0dd", 
X"a0e5", X"a0ee", X"a0f6", X"a0fe", X"a107", X"a10f", X"a118", X"a120", 
X"a129", X"a131", X"a139", X"a142", X"a14a", X"a153", X"a15b", X"a164", 
X"a16c", X"a175", X"a17d", X"a186", X"a18e", X"a197", X"a19f", X"a1a8", 
X"a1b0", X"a1b8", X"a1c1", X"a1c9", X"a1d2", X"a1db", X"a1e3", X"a1ec", 
X"a1f4", X"a1fd", X"a205", X"a20e", X"a216", X"a21f", X"a227", X"a230", 
X"a238", X"a241", X"a249", X"a252", X"a25b", X"a263", X"a26c", X"a274", 
X"a27d", X"a286", X"a28e", X"a297", X"a29f", X"a2a8", X"a2b0", X"a2b9", 
X"a2c2", X"a2ca", X"a2d3", X"a2dc", X"a2e4", X"a2ed", X"a2f5", X"a2fe", 
X"a307", X"a30f", X"a318", X"a321", X"a329", X"a332", X"a33b", X"a343", 
X"a34c", X"a355", X"a35d", X"a366", X"a36f", X"a377", X"a380", X"a389", 
X"a391", X"a39a", X"a3a3", X"a3ab", X"a3b4", X"a3bd", X"a3c6", X"a3ce", 
X"a3d7", X"a3e0", X"a3e8", X"a3f1", X"a3fa", X"a403", X"a40b", X"a414", 
X"a41d", X"a426", X"a42e", X"a437", X"a440", X"a449", X"a451", X"a45a", 
X"a463", X"a46c", X"a474", X"a47d", X"a486", X"a48f", X"a498", X"a4a0", 
X"a4a9", X"a4b2", X"a4bb", X"a4c4", X"a4cc", X"a4d5", X"a4de", X"a4e7", 
X"a4f0", X"a4f9", X"a501", X"a50a", X"a513", X"a51c", X"a525", X"a52e", 
X"a537", X"a53f", X"a548", X"a551", X"a55a", X"a563", X"a56c", X"a575", 
X"a57e", X"a586", X"a58f", X"a598", X"a5a1", X"a5aa", X"a5b3", X"a5bc", 
X"a5c5", X"a5ce", X"a5d7", X"a5df", X"a5e8", X"a5f1", X"a5fa", X"a603", 
X"a60c", X"a615", X"a61e", X"a627", X"a630", X"a639", X"a642", X"a64b", 
X"a654", X"a65d", X"a666", X"a66f", X"a678", X"a681", X"a68a", X"a693", 
X"a69c", X"a6a5", X"a6ae", X"a6b7", X"a6c0", X"a6c9", X"a6d2", X"a6db", 
X"a6e4", X"a6ed", X"a6f6", X"a6ff", X"a708", X"a711", X"a71a", X"a723", 
X"a72c", X"a735", X"a73e", X"a747", X"a750", X"a759", X"a762", X"a76b", 
X"a774", X"a77e", X"a787", X"a790", X"a799", X"a7a2", X"a7ab", X"a7b4", 
X"a7bd", X"a7c6", X"a7cf", X"a7d8", X"a7e2", X"a7eb", X"a7f4", X"a7fd", 
X"a806", X"a80f", X"a818", X"a821", X"a82b", X"a834", X"a83d", X"a846", 
X"a84f", X"a858", X"a861", X"a86b", X"a874", X"a87d", X"a886", X"a88f", 
X"a899", X"a8a2", X"a8ab", X"a8b4", X"a8bd", X"a8c6", X"a8d0", X"a8d9", 
X"a8e2", X"a8eb", X"a8f4", X"a8fe", X"a907", X"a910", X"a919", X"a923", 
X"a92c", X"a935", X"a93e", X"a948", X"a951", X"a95a", X"a963", X"a96d", 
X"a976", X"a97f", X"a988", X"a992", X"a99b", X"a9a4", X"a9ad", X"a9b7", 
X"a9c0", X"a9c9", X"a9d3", X"a9dc", X"a9e5", X"a9ee", X"a9f8", X"aa01", 
X"aa0a", X"aa14", X"aa1d", X"aa26", X"aa30", X"aa39", X"aa42", X"aa4c", 
X"aa55", X"aa5e", X"aa68", X"aa71", X"aa7a", X"aa84", X"aa8d", X"aa96", 
X"aaa0", X"aaa9", X"aab2", X"aabc", X"aac5", X"aacf", X"aad8", X"aae1", 
X"aaeb", X"aaf4", X"aafe", X"ab07", X"ab10", X"ab1a", X"ab23", X"ab2d", 
X"ab36", X"ab3f", X"ab49", X"ab52", X"ab5c", X"ab65", X"ab6f", X"ab78", 
X"ab81", X"ab8b", X"ab94", X"ab9e", X"aba7", X"abb1", X"abba", X"abc4", 
X"abcd", X"abd6", X"abe0", X"abe9", X"abf3", X"abfc", X"ac06", X"ac0f", 
X"ac19", X"ac22", X"ac2c", X"ac35", X"ac3f", X"ac48", X"ac52", X"ac5b", 
X"ac65", X"ac6e", X"ac78", X"ac81", X"ac8b", X"ac94", X"ac9e", X"aca8", 
X"acb1", X"acbb", X"acc4", X"acce", X"acd7", X"ace1", X"acea", X"acf4", 
X"acfd", X"ad07", X"ad11", X"ad1a", X"ad24", X"ad2d", X"ad37", X"ad41", 
X"ad4a", X"ad54", X"ad5d", X"ad67", X"ad70", X"ad7a", X"ad84", X"ad8d", 
X"ad97", X"ada1", X"adaa", X"adb4", X"adbd", X"adc7", X"add1", X"adda", 
X"ade4", X"adee", X"adf7", X"ae01", X"ae0b", X"ae14", X"ae1e", X"ae28", 
X"ae31", X"ae3b", X"ae45", X"ae4e", X"ae58", X"ae62", X"ae6b", X"ae75", 
X"ae7f", X"ae88", X"ae92", X"ae9c", X"aea5", X"aeaf", X"aeb9", X"aec2", 
X"aecc", X"aed6", X"aee0", X"aee9", X"aef3", X"aefd", X"af07", X"af10", 
X"af1a", X"af24", X"af2d", X"af37", X"af41", X"af4b", X"af54", X"af5e", 
X"af68", X"af72", X"af7c", X"af85", X"af8f", X"af99", X"afa3", X"afac", 
X"afb6", X"afc0", X"afca", X"afd4", X"afdd", X"afe7", X"aff1", X"affb", 
X"b005", X"b00e", X"b018", X"b022", X"b02c", X"b036", X"b040", X"b049", 
X"b053", X"b05d", X"b067", X"b071", X"b07b", X"b084", X"b08e", X"b098", 
X"b0a2", X"b0ac", X"b0b6", X"b0c0", X"b0c9", X"b0d3", X"b0dd", X"b0e7", 
X"b0f1", X"b0fb", X"b105", X"b10f", X"b118", X"b122", X"b12c", X"b136", 
X"b140", X"b14a", X"b154", X"b15e", X"b168", X"b172", X"b17c", X"b186", 
X"b18f", X"b199", X"b1a3", X"b1ad", X"b1b7", X"b1c1", X"b1cb", X"b1d5", 
X"b1df", X"b1e9", X"b1f3", X"b1fd", X"b207", X"b211", X"b21b", X"b225", 
X"b22f", X"b239", X"b243", X"b24d", X"b257", X"b261", X"b26b", X"b275", 
X"b27f", X"b289", X"b293", X"b29d", X"b2a7", X"b2b1", X"b2bb", X"b2c5", 
X"b2cf", X"b2d9", X"b2e3", X"b2ed", X"b2f7", X"b301", X"b30b", X"b315", 
X"b31f", X"b329", X"b333", X"b33d", X"b347", X"b351", X"b35b", X"b365", 
X"b36f", X"b37a", X"b384", X"b38e", X"b398", X"b3a2", X"b3ac", X"b3b6", 
X"b3c0", X"b3ca", X"b3d4", X"b3de", X"b3e9", X"b3f3", X"b3fd", X"b407", 
X"b411", X"b41b", X"b425", X"b42f", X"b439", X"b444", X"b44e", X"b458", 
X"b462", X"b46c", X"b476", X"b480", X"b48b", X"b495", X"b49f", X"b4a9", 
X"b4b3", X"b4bd", X"b4c8", X"b4d2", X"b4dc", X"b4e6", X"b4f0", X"b4fa", 
X"b505", X"b50f", X"b519", X"b523", X"b52d", X"b538", X"b542", X"b54c", 
X"b556", X"b560", X"b56b", X"b575", X"b57f", X"b589", X"b593", X"b59e", 
X"b5a8", X"b5b2", X"b5bc", X"b5c7", X"b5d1", X"b5db", X"b5e5", X"b5f0", 
X"b5fa", X"b604", X"b60e", X"b619", X"b623", X"b62d", X"b637", X"b642", 
X"b64c", X"b656", X"b660", X"b66b", X"b675", X"b67f", X"b68a", X"b694", 
X"b69e", X"b6a8", X"b6b3", X"b6bd", X"b6c7", X"b6d2", X"b6dc", X"b6e6", 
X"b6f1", X"b6fb", X"b705", X"b710", X"b71a", X"b724", X"b72f", X"b739", 
X"b743", X"b74e", X"b758", X"b762", X"b76d", X"b777", X"b781", X"b78c", 
X"b796", X"b7a0", X"b7ab", X"b7b5", X"b7c0", X"b7ca", X"b7d4", X"b7df", 
X"b7e9", X"b7f3", X"b7fe", X"b808", X"b813", X"b81d", X"b827", X"b832", 
X"b83c", X"b847", X"b851", X"b85b", X"b866", X"b870", X"b87b", X"b885", 
X"b890", X"b89a", X"b8a4", X"b8af", X"b8b9", X"b8c4", X"b8ce", X"b8d9", 
X"b8e3", X"b8ee", X"b8f8", X"b902", X"b90d", X"b917", X"b922", X"b92c", 
X"b937", X"b941", X"b94c", X"b956", X"b961", X"b96b", X"b976", X"b980", 
X"b98b", X"b995", X"b9a0", X"b9aa", X"b9b5", X"b9bf", X"b9ca", X"b9d4", 
X"b9df", X"b9e9", X"b9f4", X"b9fe", X"ba09", X"ba13", X"ba1e", X"ba28", 
X"ba33", X"ba3d", X"ba48", X"ba52", X"ba5d", X"ba67", X"ba72", X"ba7d", 
X"ba87", X"ba92", X"ba9c", X"baa7", X"bab1", X"babc", X"bac7", X"bad1", 
X"badc", X"bae6", X"baf1", X"bafb", X"bb06", X"bb11", X"bb1b", X"bb26", 
X"bb30", X"bb3b", X"bb46", X"bb50", X"bb5b", X"bb65", X"bb70", X"bb7b", 
X"bb85", X"bb90", X"bb9a", X"bba5", X"bbb0", X"bbba", X"bbc5", X"bbd0", 
X"bbda", X"bbe5", X"bbef", X"bbfa", X"bc05", X"bc0f", X"bc1a", X"bc25", 
X"bc2f", X"bc3a", X"bc45", X"bc4f", X"bc5a", X"bc65", X"bc6f", X"bc7a", 
X"bc85", X"bc8f", X"bc9a", X"bca5", X"bcaf", X"bcba", X"bcc5", X"bcd0", 
X"bcda", X"bce5", X"bcf0", X"bcfa", X"bd05", X"bd10", X"bd1a", X"bd25", 
X"bd30", X"bd3b", X"bd45", X"bd50", X"bd5b", X"bd66", X"bd70", X"bd7b", 
X"bd86", X"bd90", X"bd9b", X"bda6", X"bdb1", X"bdbb", X"bdc6", X"bdd1", 
X"bddc", X"bde6", X"bdf1", X"bdfc", X"be07", X"be12", X"be1c", X"be27", 
X"be32", X"be3d", X"be47", X"be52", X"be5d", X"be68", X"be73", X"be7d", 
X"be88", X"be93", X"be9e", X"bea9", X"beb3", X"bebe", X"bec9", X"bed4", 
X"bedf", X"bee9", X"bef4", X"beff", X"bf0a", X"bf15", X"bf20", X"bf2a", 
X"bf35", X"bf40", X"bf4b", X"bf56", X"bf61", X"bf6b", X"bf76", X"bf81", 
X"bf8c", X"bf97", X"bfa2", X"bfad", X"bfb8", X"bfc2", X"bfcd", X"bfd8", 
X"bfe3", X"bfee", X"bff9", X"c004", X"c00f", X"c019", X"c024", X"c02f", 
X"c03a", X"c045", X"c050", X"c05b", X"c066", X"c071", X"c07b", X"c086", 
X"c091", X"c09c", X"c0a7", X"c0b2", X"c0bd", X"c0c8", X"c0d3", X"c0de", 
X"c0e9", X"c0f4", X"c0ff", X"c10a", X"c114", X"c11f", X"c12a", X"c135", 
X"c140", X"c14b", X"c156", X"c161", X"c16c", X"c177", X"c182", X"c18d", 
X"c198", X"c1a3", X"c1ae", X"c1b9", X"c1c4", X"c1cf", X"c1da", X"c1e5", 
X"c1f0", X"c1fb", X"c206", X"c211", X"c21c", X"c227", X"c232", X"c23d", 
X"c248", X"c253", X"c25e", X"c269", X"c274", X"c27f", X"c28a", X"c295", 
X"c2a0", X"c2ab", X"c2b6", X"c2c1", X"c2cc", X"c2d7", X"c2e2", X"c2ed", 
X"c2f8", X"c303", X"c30e", X"c319", X"c324", X"c330", X"c33b", X"c346", 
X"c351", X"c35c", X"c367", X"c372", X"c37d", X"c388", X"c393", X"c39e", 
X"c3a9", X"c3b4", X"c3bf", X"c3cb", X"c3d6", X"c3e1", X"c3ec", X"c3f7", 
X"c402", X"c40d", X"c418", X"c423", X"c42e", X"c43a", X"c445", X"c450", 
X"c45b", X"c466", X"c471", X"c47c", X"c487", X"c493", X"c49e", X"c4a9", 
X"c4b4", X"c4bf", X"c4ca", X"c4d5", X"c4e0", X"c4ec", X"c4f7", X"c502", 
X"c50d", X"c518", X"c523", X"c52f", X"c53a", X"c545", X"c550", X"c55b", 
X"c566", X"c572", X"c57d", X"c588", X"c593", X"c59e", X"c5a9", X"c5b5", 
X"c5c0", X"c5cb", X"c5d6", X"c5e1", X"c5ed", X"c5f8", X"c603", X"c60e", 
X"c619", X"c625", X"c630", X"c63b", X"c646", X"c651", X"c65d", X"c668", 
X"c673", X"c67e", X"c68a", X"c695", X"c6a0", X"c6ab", X"c6b7", X"c6c2", 
X"c6cd", X"c6d8", X"c6e3", X"c6ef", X"c6fa", X"c705", X"c710", X"c71c", 
X"c727", X"c732", X"c73e", X"c749", X"c754", X"c75f", X"c76b", X"c776", 
X"c781", X"c78c", X"c798", X"c7a3", X"c7ae", X"c7ba", X"c7c5", X"c7d0", 
X"c7db", X"c7e7", X"c7f2", X"c7fd", X"c809", X"c814", X"c81f", X"c82b", 
X"c836", X"c841", X"c84c", X"c858", X"c863", X"c86e", X"c87a", X"c885", 
X"c890", X"c89c", X"c8a7", X"c8b2", X"c8be", X"c8c9", X"c8d4", X"c8e0", 
X"c8eb", X"c8f6", X"c902", X"c90d", X"c918", X"c924", X"c92f", X"c93b", 
X"c946", X"c951", X"c95d", X"c968", X"c973", X"c97f", X"c98a", X"c995", 
X"c9a1", X"c9ac", X"c9b8", X"c9c3", X"c9ce", X"c9da", X"c9e5", X"c9f1", 
X"c9fc", X"ca07", X"ca13", X"ca1e", X"ca29", X"ca35", X"ca40", X"ca4c", 
X"ca57", X"ca63", X"ca6e", X"ca79", X"ca85", X"ca90", X"ca9c", X"caa7", 
X"cab2", X"cabe", X"cac9", X"cad5", X"cae0", X"caec", X"caf7", X"cb02", 
X"cb0e", X"cb19", X"cb25", X"cb30", X"cb3c", X"cb47", X"cb53", X"cb5e", 
X"cb69", X"cb75", X"cb80", X"cb8c", X"cb97", X"cba3", X"cbae", X"cbba", 
X"cbc5", X"cbd1", X"cbdc", X"cbe8", X"cbf3", X"cbff", X"cc0a", X"cc16", 
X"cc21", X"cc2d", X"cc38", X"cc44", X"cc4f", X"cc5b", X"cc66", X"cc72", 
X"cc7d", X"cc89", X"cc94", X"cca0", X"ccab", X"ccb7", X"ccc2", X"ccce", 
X"ccd9", X"cce5", X"ccf0", X"ccfc", X"cd07", X"cd13", X"cd1e", X"cd2a", 
X"cd35", X"cd41", X"cd4c", X"cd58", X"cd63", X"cd6f", X"cd7b", X"cd86", 
X"cd92", X"cd9d", X"cda9", X"cdb4", X"cdc0", X"cdcb", X"cdd7", X"cde3", 
X"cdee", X"cdfa", X"ce05", X"ce11", X"ce1c", X"ce28", X"ce34", X"ce3f", 
X"ce4b", X"ce56", X"ce62", X"ce6d", X"ce79", X"ce85", X"ce90", X"ce9c", 
X"cea7", X"ceb3", X"cebf", X"ceca", X"ced6", X"cee1", X"ceed", X"cef9", 
X"cf04", X"cf10", X"cf1b", X"cf27", X"cf33", X"cf3e", X"cf4a", X"cf56", 
X"cf61", X"cf6d", X"cf78", X"cf84", X"cf90", X"cf9b", X"cfa7", X"cfb3", 
X"cfbe", X"cfca", X"cfd6", X"cfe1", X"cfed", X"cff8", X"d004", X"d010", 
X"d01b", X"d027", X"d033", X"d03e", X"d04a", X"d056", X"d061", X"d06d", 
X"d079", X"d084", X"d090", X"d09c", X"d0a7", X"d0b3", X"d0bf", X"d0ca", 
X"d0d6", X"d0e2", X"d0ed", X"d0f9", X"d105", X"d111", X"d11c", X"d128", 
X"d134", X"d13f", X"d14b", X"d157", X"d162", X"d16e", X"d17a", X"d186", 
X"d191", X"d19d", X"d1a9", X"d1b4", X"d1c0", X"d1cc", X"d1d8", X"d1e3", 
X"d1ef", X"d1fb", X"d206", X"d212", X"d21e", X"d22a", X"d235", X"d241", 
X"d24d", X"d259", X"d264", X"d270", X"d27c", X"d288", X"d293", X"d29f", 
X"d2ab", X"d2b7", X"d2c2", X"d2ce", X"d2da", X"d2e6", X"d2f1", X"d2fd", 
X"d309", X"d315", X"d320", X"d32c", X"d338", X"d344", X"d34f", X"d35b", 
X"d367", X"d373", X"d37f", X"d38a", X"d396", X"d3a2", X"d3ae", X"d3ba", 
X"d3c5", X"d3d1", X"d3dd", X"d3e9", X"d3f4", X"d400", X"d40c", X"d418", 
X"d424", X"d430", X"d43b", X"d447", X"d453", X"d45f", X"d46b", X"d476", 
X"d482", X"d48e", X"d49a", X"d4a6", X"d4b1", X"d4bd", X"d4c9", X"d4d5", 
X"d4e1", X"d4ed", X"d4f8", X"d504", X"d510", X"d51c", X"d528", X"d534", 
X"d53f", X"d54b", X"d557", X"d563", X"d56f", X"d57b", X"d587", X"d592", 
X"d59e", X"d5aa", X"d5b6", X"d5c2", X"d5ce", X"d5da", X"d5e5", X"d5f1", 
X"d5fd", X"d609", X"d615", X"d621", X"d62d", X"d639", X"d644", X"d650", 
X"d65c", X"d668", X"d674", X"d680", X"d68c", X"d698", X"d6a4", X"d6af", 
X"d6bb", X"d6c7", X"d6d3", X"d6df", X"d6eb", X"d6f7", X"d703", X"d70f", 
X"d71b", X"d726", X"d732", X"d73e", X"d74a", X"d756", X"d762", X"d76e", 
X"d77a", X"d786", X"d792", X"d79e", X"d7aa", X"d7b5", X"d7c1", X"d7cd", 
X"d7d9", X"d7e5", X"d7f1", X"d7fd", X"d809", X"d815", X"d821", X"d82d", 
X"d839", X"d845", X"d851", X"d85d", X"d869", X"d875", X"d880", X"d88c", 
X"d898", X"d8a4", X"d8b0", X"d8bc", X"d8c8", X"d8d4", X"d8e0", X"d8ec", 
X"d8f8", X"d904", X"d910", X"d91c", X"d928", X"d934", X"d940", X"d94c", 
X"d958", X"d964", X"d970", X"d97c", X"d988", X"d994", X"d9a0", X"d9ac", 
X"d9b8", X"d9c4", X"d9d0", X"d9dc", X"d9e8", X"d9f4", X"da00", X"da0c", 
X"da18", X"da24", X"da30", X"da3c", X"da48", X"da54", X"da60", X"da6c", 
X"da78", X"da84", X"da90", X"da9c", X"daa8", X"dab4", X"dac0", X"dacc", 
X"dad8", X"dae4", X"daf0", X"dafc", X"db08", X"db14", X"db20", X"db2c", 
X"db38", X"db44", X"db50", X"db5c", X"db68", X"db74", X"db80", X"db8c", 
X"db99", X"dba5", X"dbb1", X"dbbd", X"dbc9", X"dbd5", X"dbe1", X"dbed", 
X"dbf9", X"dc05", X"dc11", X"dc1d", X"dc29", X"dc35", X"dc41", X"dc4d", 
X"dc59", X"dc66", X"dc72", X"dc7e", X"dc8a", X"dc96", X"dca2", X"dcae", 
X"dcba", X"dcc6", X"dcd2", X"dcde", X"dcea", X"dcf6", X"dd03", X"dd0f", 
X"dd1b", X"dd27", X"dd33", X"dd3f", X"dd4b", X"dd57", X"dd63", X"dd6f", 
X"dd7c", X"dd88", X"dd94", X"dda0", X"ddac", X"ddb8", X"ddc4", X"ddd0", 
X"dddc", X"dde8", X"ddf5", X"de01", X"de0d", X"de19", X"de25", X"de31", 
X"de3d", X"de49", X"de56", X"de62", X"de6e", X"de7a", X"de86", X"de92", 
X"de9e", X"deaa", X"deb7", X"dec3", X"decf", X"dedb", X"dee7", X"def3", 
X"deff", X"df0c", X"df18", X"df24", X"df30", X"df3c", X"df48", X"df54", 
X"df61", X"df6d", X"df79", X"df85", X"df91", X"df9d", X"dfa9", X"dfb6", 
X"dfc2", X"dfce", X"dfda", X"dfe6", X"dff2", X"dfff", X"e00b", X"e017", 
X"e023", X"e02f", X"e03b", X"e048", X"e054", X"e060", X"e06c", X"e078", 
X"e085", X"e091", X"e09d", X"e0a9", X"e0b5", X"e0c1", X"e0ce", X"e0da", 
X"e0e6", X"e0f2", X"e0fe", X"e10b", X"e117", X"e123", X"e12f", X"e13b", 
X"e148", X"e154", X"e160", X"e16c", X"e178", X"e185", X"e191", X"e19d", 
X"e1a9", X"e1b5", X"e1c2", X"e1ce", X"e1da", X"e1e6", X"e1f2", X"e1ff", 
X"e20b", X"e217", X"e223", X"e230", X"e23c", X"e248", X"e254", X"e260", 
X"e26d", X"e279", X"e285", X"e291", X"e29e", X"e2aa", X"e2b6", X"e2c2", 
X"e2cf", X"e2db", X"e2e7", X"e2f3", X"e2ff", X"e30c", X"e318", X"e324", 
X"e330", X"e33d", X"e349", X"e355", X"e361", X"e36e", X"e37a", X"e386", 
X"e392", X"e39f", X"e3ab", X"e3b7", X"e3c3", X"e3d0", X"e3dc", X"e3e8", 
X"e3f4", X"e401", X"e40d", X"e419", X"e426", X"e432", X"e43e", X"e44a", 
X"e457", X"e463", X"e46f", X"e47b", X"e488", X"e494", X"e4a0", X"e4ad", 
X"e4b9", X"e4c5", X"e4d1", X"e4de", X"e4ea", X"e4f6", X"e502", X"e50f", 
X"e51b", X"e527", X"e534", X"e540", X"e54c", X"e558", X"e565", X"e571", 
X"e57d", X"e58a", X"e596", X"e5a2", X"e5af", X"e5bb", X"e5c7", X"e5d3", 
X"e5e0", X"e5ec", X"e5f8", X"e605", X"e611", X"e61d", X"e62a", X"e636", 
X"e642", X"e64f", X"e65b", X"e667", X"e673", X"e680", X"e68c", X"e698", 
X"e6a5", X"e6b1", X"e6bd", X"e6ca", X"e6d6", X"e6e2", X"e6ef", X"e6fb", 
X"e707", X"e714", X"e720", X"e72c", X"e739", X"e745", X"e751", X"e75e", 
X"e76a", X"e776", X"e783", X"e78f", X"e79b", X"e7a8", X"e7b4", X"e7c0", 
X"e7cd", X"e7d9", X"e7e5", X"e7f2", X"e7fe", X"e80a", X"e817", X"e823", 
X"e82f", X"e83c", X"e848", X"e854", X"e861", X"e86d", X"e879", X"e886", 
X"e892", X"e89f", X"e8ab", X"e8b7", X"e8c4", X"e8d0", X"e8dc", X"e8e9", 
X"e8f5", X"e901", X"e90e", X"e91a", X"e926", X"e933", X"e93f", X"e94c", 
X"e958", X"e964", X"e971", X"e97d", X"e989", X"e996", X"e9a2", X"e9af", 
X"e9bb", X"e9c7", X"e9d4", X"e9e0", X"e9ec", X"e9f9", X"ea05", X"ea12", 
X"ea1e", X"ea2a", X"ea37", X"ea43", X"ea4f", X"ea5c", X"ea68", X"ea75", 
X"ea81", X"ea8d", X"ea9a", X"eaa6", X"eab3", X"eabf", X"eacb", X"ead8", 
X"eae4", X"eaf1", X"eafd", X"eb09", X"eb16", X"eb22", X"eb2f", X"eb3b", 
X"eb47", X"eb54", X"eb60", X"eb6d", X"eb79", X"eb85", X"eb92", X"eb9e", 
X"ebab", X"ebb7", X"ebc3", X"ebd0", X"ebdc", X"ebe9", X"ebf5", X"ec01", 
X"ec0e", X"ec1a", X"ec27", X"ec33", X"ec3f", X"ec4c", X"ec58", X"ec65", 
X"ec71", X"ec7e", X"ec8a", X"ec96", X"eca3", X"ecaf", X"ecbc", X"ecc8", 
X"ecd5", X"ece1", X"eced", X"ecfa", X"ed06", X"ed13", X"ed1f", X"ed2c", 
X"ed38", X"ed44", X"ed51", X"ed5d", X"ed6a", X"ed76", X"ed83", X"ed8f", 
X"ed9b", X"eda8", X"edb4", X"edc1", X"edcd", X"edda", X"ede6", X"edf2", 
X"edff", X"ee0b", X"ee18", X"ee24", X"ee31", X"ee3d", X"ee4a", X"ee56", 
X"ee62", X"ee6f", X"ee7b", X"ee88", X"ee94", X"eea1", X"eead", X"eeba", 
X"eec6", X"eed3", X"eedf", X"eeeb", X"eef8", X"ef04", X"ef11", X"ef1d", 
X"ef2a", X"ef36", X"ef43", X"ef4f", X"ef5c", X"ef68", X"ef74", X"ef81", 
X"ef8d", X"ef9a", X"efa6", X"efb3", X"efbf", X"efcc", X"efd8", X"efe5", 
X"eff1", X"effe", X"f00a", X"f016", X"f023", X"f02f", X"f03c", X"f048", 
X"f055", X"f061", X"f06e", X"f07a", X"f087", X"f093", X"f0a0", X"f0ac", 
X"f0b9", X"f0c5", X"f0d2", X"f0de", X"f0eb", X"f0f7", X"f104", X"f110", 
X"f11c", X"f129", X"f135", X"f142", X"f14e", X"f15b", X"f167", X"f174", 
X"f180", X"f18d", X"f199", X"f1a6", X"f1b2", X"f1bf", X"f1cb", X"f1d8", 
X"f1e4", X"f1f1", X"f1fd", X"f20a", X"f216", X"f223", X"f22f", X"f23c", 
X"f248", X"f255", X"f261", X"f26e", X"f27a", X"f287", X"f293", X"f2a0", 
X"f2ac", X"f2b9", X"f2c5", X"f2d2", X"f2de", X"f2eb", X"f2f7", X"f304", 
X"f310", X"f31d", X"f329", X"f336", X"f342", X"f34f", X"f35b", X"f368", 
X"f374", X"f381", X"f38d", X"f39a", X"f3a6", X"f3b3", X"f3bf", X"f3cc", 
X"f3d8", X"f3e5", X"f3f1", X"f3fe", X"f40a", X"f417", X"f423", X"f430", 
X"f43c", X"f449", X"f455", X"f462", X"f46e", X"f47b", X"f487", X"f494", 
X"f4a0", X"f4ad", X"f4b9", X"f4c6", X"f4d3", X"f4df", X"f4ec", X"f4f8", 
X"f505", X"f511", X"f51e", X"f52a", X"f537", X"f543", X"f550", X"f55c", 
X"f569", X"f575", X"f582", X"f58e", X"f59b", X"f5a7", X"f5b4", X"f5c0", 
X"f5cd", X"f5d9", X"f5e6", X"f5f3", X"f5ff", X"f60c", X"f618", X"f625", 
X"f631", X"f63e", X"f64a", X"f657", X"f663", X"f670", X"f67c", X"f689", 
X"f695", X"f6a2", X"f6af", X"f6bb", X"f6c8", X"f6d4", X"f6e1", X"f6ed", 
X"f6fa", X"f706", X"f713", X"f71f", X"f72c", X"f738", X"f745", X"f751", 
X"f75e", X"f76b", X"f777", X"f784", X"f790", X"f79d", X"f7a9", X"f7b6", 
X"f7c2", X"f7cf", X"f7db", X"f7e8", X"f7f4", X"f801", X"f80e", X"f81a", 
X"f827", X"f833", X"f840", X"f84c", X"f859", X"f865", X"f872", X"f87e", 
X"f88b", X"f898", X"f8a4", X"f8b1", X"f8bd", X"f8ca", X"f8d6", X"f8e3", 
X"f8ef", X"f8fc", X"f908", X"f915", X"f922", X"f92e", X"f93b", X"f947", 
X"f954", X"f960", X"f96d", X"f979", X"f986", X"f992", X"f99f", X"f9ac", 
X"f9b8", X"f9c5", X"f9d1", X"f9de", X"f9ea", X"f9f7", X"fa03", X"fa10", 
X"fa1d", X"fa29", X"fa36", X"fa42", X"fa4f", X"fa5b", X"fa68", X"fa74", 
X"fa81", X"fa8e", X"fa9a", X"faa7", X"fab3", X"fac0", X"facc", X"fad9", 
X"fae5", X"faf2", X"faff", X"fb0b", X"fb18", X"fb24", X"fb31", X"fb3d", 
X"fb4a", X"fb56", X"fb63", X"fb70", X"fb7c", X"fb89", X"fb95", X"fba2", 
X"fbae", X"fbbb", X"fbc7", X"fbd4", X"fbe1", X"fbed", X"fbfa", X"fc06", 
X"fc13", X"fc1f", X"fc2c", X"fc39", X"fc45", X"fc52", X"fc5e", X"fc6b", 
X"fc77", X"fc84", X"fc90", X"fc9d", X"fcaa", X"fcb6", X"fcc3", X"fccf", 
X"fcdc", X"fce8", X"fcf5", X"fd02", X"fd0e", X"fd1b", X"fd27", X"fd34", 
X"fd40", X"fd4d", X"fd59", X"fd66", X"fd73", X"fd7f", X"fd8c", X"fd98", 
X"fda5", X"fdb1", X"fdbe", X"fdcb", X"fdd7", X"fde4", X"fdf0", X"fdfd", 
X"fe09", X"fe16", X"fe22", X"fe2f", X"fe3c", X"fe48", X"fe55", X"fe61", 
X"fe6e", X"fe7a", X"fe87", X"fe94", X"fea0", X"fead", X"feb9", X"fec6", 
X"fed2", X"fedf", X"feec", X"fef8", X"ff05", X"ff11", X"ff1e", X"ff2a", 
X"ff37", X"ff44", X"ff50", X"ff5d", X"ff69", X"ff76", X"ff82", X"ff8f", 
X"ff9b", X"ffa8", X"ffb5", X"ffc1", X"ffce", X"ffda", X"ffe7", X"fff3" 
);

signal counter : std_logic := '0';
signal value : std_logic_vector(15 downto 0);
signal current_addr:std_logic_vector(13 downto 0);
begin

rom_select: process (clk)
begin
  if rising_edge(clk) then
	 counter <= not counter;
    value <= SIN_ROM(conv_integer(current_addr)) + 8192;
	 if counter = '0' then
      current_addr <= addr;
		sin_out <= value;
	 else
      current_addr <= addr_1;
		sin_out_1 <= value;
	  end if;
	
  end if;
end process rom_select;


end rtl;